magic
tech sky130A
magscale 1 2
timestamp 1712843699
<< metal1 >>
rect -900 10600 -700 10820
rect -900 10480 -860 10600
rect -740 10480 -700 10600
rect -900 10440 -700 10480
rect 700 3920 1160 4040
rect 580 3740 1280 3920
rect 580 3720 2400 3740
rect -320 3560 -160 3580
rect -320 3440 -300 3560
rect -180 3440 -160 3560
rect -320 2640 -160 3440
rect 580 3560 2220 3720
rect 2380 3560 2400 3720
rect 8000 3700 8200 3740
rect 7740 3680 8200 3700
rect 7740 3580 7760 3680
rect 7880 3580 8200 3680
rect 7740 3560 8200 3580
rect 580 3540 2400 3560
rect 8000 3540 8200 3560
rect 580 3140 1280 3540
rect -400 2440 1280 2640
rect -540 2320 -80 2440
rect -660 1560 40 2320
rect 640 2120 1220 2180
rect -540 740 280 940
rect -620 520 -20 580
rect 80 380 280 740
rect -900 360 1800 380
rect -900 200 1620 360
rect 1780 200 1800 360
rect -900 180 1800 200
<< via1 >>
rect -860 10480 -740 10600
rect -300 3440 -180 3560
rect 2220 3560 2380 3720
rect 7760 3580 7880 3680
rect 1620 200 1780 360
<< metal2 >>
rect -860 10600 -740 10610
rect -860 10470 -740 10480
rect 2220 3720 2380 3730
rect -300 3560 -180 3570
rect 7760 3680 7880 3690
rect 7760 3570 7880 3580
rect 2220 3550 2380 3560
rect -300 3430 -180 3440
rect 1620 360 1780 370
rect 1620 190 1780 200
<< via2 >>
rect -860 10480 -740 10600
rect -300 3440 -180 3560
rect 2220 3560 2380 3720
rect 7760 3580 7880 3680
rect 1620 200 1780 360
<< metal3 >>
rect -870 10600 -730 10605
rect -870 10480 -860 10600
rect -740 10480 -730 10600
rect -870 10475 -730 10480
rect 2210 3720 2390 3725
rect -310 3560 -170 3565
rect -310 3440 -300 3560
rect -180 3440 -170 3560
rect 2210 3560 2220 3720
rect 2380 3560 2390 3720
rect 7750 3680 7890 3685
rect 7750 3580 7760 3680
rect 7880 3580 7890 3680
rect 7750 3575 7890 3580
rect 2210 3555 2390 3560
rect -310 3435 -170 3440
rect 1790 365 1800 385
rect 1610 360 1800 365
rect 1610 200 1620 360
rect 1780 200 1800 360
rect 1610 195 1800 200
rect 1790 175 1800 195
<< via3 >>
rect -860 10480 -740 10600
rect -300 3440 -180 3560
rect 2220 3560 2380 3720
rect 7760 3580 7880 3680
rect 1620 200 1780 360
<< metal4 >>
rect -861 10600 -739 10601
rect -861 10480 -860 10600
rect -740 10480 -739 10600
rect -861 10479 -739 10480
rect -840 10380 -740 10479
rect -840 10280 -700 10380
rect -800 10220 -700 10280
rect -320 3560 -160 4360
rect -320 3440 -300 3560
rect -180 3440 -160 3560
rect -320 3420 -160 3440
rect 2200 3720 2400 3740
rect 2200 3560 2220 3720
rect 2380 3560 2400 3720
rect 2200 3280 2400 3560
rect 7740 3680 7900 3700
rect 7740 3580 7760 3680
rect 7880 3580 7900 3680
rect 7740 3280 7900 3580
rect 1600 360 1880 380
rect 1600 200 1620 360
rect 1780 200 1880 360
rect 1600 180 1880 200
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1712795588
transform -1 0 2349 0 1 7180
box -3150 -3100 3149 3100
use sky130_fd_pr__cap_mim_m3_1_3MBNLG  XC3
timestamp 1712843110
transform -1 0 4949 0 1 -5950
box -3150 -9450 3149 9450
use sky130_fd_pr__pfet_01v8_lvt_3F9YD3  sky130_fd_pr__pfet_01v8_lvt_3F9YD3_0
timestamp 1712834386
transform 1 0 -313 0 1 1419
box -487 -1019 487 1019
use sky130_fd_pr__pfet_01v8_lvt_3F9YD3  sky130_fd_pr__pfet_01v8_lvt_3F9YD3_1
timestamp 1712834386
transform 1 0 927 0 1 3019
box -487 -1019 487 1019
<< labels >>
flabel metal1 -900 180 -700 380 0 FreeSans 256 0 0 0 ground
port 0 nsew
flabel metal1 -900 10620 -700 10820 0 FreeSans 256 0 0 0 i
port 2 nsew
flabel metal1 8000 3540 8200 3740 0 FreeSans 256 0 0 0 o
port 1 nsew
<< end >>
