magic
tech sky130A
magscale 1 2
timestamp 1712949221
<< nwell >>
rect 1100 22900 2074 24938
rect 2340 24500 3314 26538
rect 10240 22900 11214 24938
rect 11480 24500 12454 26538
rect 19430 22900 20404 24938
rect 20670 24500 21644 26538
rect 28560 18140 32372 19334
rect 29850 15890 32372 18140
rect 32630 16840 33246 18754
<< pwell >>
rect 31167 25401 33683 25957
rect 30172 19392 32376 20508
rect 33302 15892 33858 19708
<< nnmos >>
rect 31425 25629 33425 25729
<< mvnmos >>
rect 30400 19650 30600 20250
rect 30658 19650 30858 20250
rect 30916 19650 31116 20250
rect 31174 19650 31374 20250
rect 31432 19650 31632 20250
rect 31690 19650 31890 20250
rect 31948 19650 32148 20250
rect 33530 18050 33630 19450
rect 33530 16150 33630 17550
<< mvpmos >>
rect 28818 18437 29018 19037
rect 29076 18437 29276 19037
rect 29334 18437 29534 19037
rect 29592 18437 29792 19037
rect 29850 18437 30050 19037
rect 30108 18437 30308 19037
rect 30366 18437 30566 19037
rect 30624 18437 30824 19037
rect 30882 18437 31082 19037
rect 31140 18437 31340 19037
rect 31398 18437 31598 19037
rect 31656 18437 31856 19037
rect 31914 18437 32114 19037
rect 30108 17317 30308 17917
rect 30366 17317 30566 17917
rect 30624 17317 30824 17917
rect 30882 17317 31082 17917
rect 31140 17317 31340 17917
rect 31398 17317 31598 17917
rect 31656 17317 31856 17917
rect 31914 17317 32114 17917
rect 32888 18057 32988 18457
rect 30108 16187 30308 16787
rect 30366 16187 30566 16787
rect 30624 16187 30824 16787
rect 30882 16187 31082 16787
rect 31140 16187 31340 16787
rect 31398 16187 31598 16787
rect 31656 16187 31856 16787
rect 31914 16187 32114 16787
rect 32888 17137 32988 17537
<< pmoslvt >>
rect 1296 23119 1366 24719
rect 1424 23119 1494 24719
rect 1552 23119 1622 24719
rect 1680 23119 1750 24719
rect 1808 23119 1878 24719
rect 2536 24719 2606 26319
rect 2664 24719 2734 26319
rect 2792 24719 2862 26319
rect 2920 24719 2990 26319
rect 3048 24719 3118 26319
rect 10436 23119 10506 24719
rect 10564 23119 10634 24719
rect 10692 23119 10762 24719
rect 10820 23119 10890 24719
rect 10948 23119 11018 24719
rect 11676 24719 11746 26319
rect 11804 24719 11874 26319
rect 11932 24719 12002 26319
rect 12060 24719 12130 26319
rect 12188 24719 12258 26319
rect 19626 23119 19696 24719
rect 19754 23119 19824 24719
rect 19882 23119 19952 24719
rect 20010 23119 20080 24719
rect 20138 23119 20208 24719
rect 20866 24719 20936 26319
rect 20994 24719 21064 26319
rect 21122 24719 21192 26319
rect 21250 24719 21320 26319
rect 21378 24719 21448 26319
<< pdiff >>
rect 1238 24707 1296 24719
rect 1238 23131 1250 24707
rect 1284 23131 1296 24707
rect 1238 23119 1296 23131
rect 1366 24707 1424 24719
rect 1366 23131 1378 24707
rect 1412 23131 1424 24707
rect 1366 23119 1424 23131
rect 1494 24707 1552 24719
rect 1494 23131 1506 24707
rect 1540 23131 1552 24707
rect 1494 23119 1552 23131
rect 1622 24707 1680 24719
rect 1622 23131 1634 24707
rect 1668 23131 1680 24707
rect 1622 23119 1680 23131
rect 1750 24707 1808 24719
rect 1750 23131 1762 24707
rect 1796 23131 1808 24707
rect 1750 23119 1808 23131
rect 1878 24707 1936 24719
rect 1878 23131 1890 24707
rect 1924 23131 1936 24707
rect 1878 23119 1936 23131
rect 2478 26307 2536 26319
rect 2478 24731 2490 26307
rect 2524 24731 2536 26307
rect 2478 24719 2536 24731
rect 2606 26307 2664 26319
rect 2606 24731 2618 26307
rect 2652 24731 2664 26307
rect 2606 24719 2664 24731
rect 2734 26307 2792 26319
rect 2734 24731 2746 26307
rect 2780 24731 2792 26307
rect 2734 24719 2792 24731
rect 2862 26307 2920 26319
rect 2862 24731 2874 26307
rect 2908 24731 2920 26307
rect 2862 24719 2920 24731
rect 2990 26307 3048 26319
rect 2990 24731 3002 26307
rect 3036 24731 3048 26307
rect 2990 24719 3048 24731
rect 3118 26307 3176 26319
rect 3118 24731 3130 26307
rect 3164 24731 3176 26307
rect 3118 24719 3176 24731
rect 10378 24707 10436 24719
rect 10378 23131 10390 24707
rect 10424 23131 10436 24707
rect 10378 23119 10436 23131
rect 10506 24707 10564 24719
rect 10506 23131 10518 24707
rect 10552 23131 10564 24707
rect 10506 23119 10564 23131
rect 10634 24707 10692 24719
rect 10634 23131 10646 24707
rect 10680 23131 10692 24707
rect 10634 23119 10692 23131
rect 10762 24707 10820 24719
rect 10762 23131 10774 24707
rect 10808 23131 10820 24707
rect 10762 23119 10820 23131
rect 10890 24707 10948 24719
rect 10890 23131 10902 24707
rect 10936 23131 10948 24707
rect 10890 23119 10948 23131
rect 11018 24707 11076 24719
rect 11018 23131 11030 24707
rect 11064 23131 11076 24707
rect 11018 23119 11076 23131
rect 11618 26307 11676 26319
rect 11618 24731 11630 26307
rect 11664 24731 11676 26307
rect 11618 24719 11676 24731
rect 11746 26307 11804 26319
rect 11746 24731 11758 26307
rect 11792 24731 11804 26307
rect 11746 24719 11804 24731
rect 11874 26307 11932 26319
rect 11874 24731 11886 26307
rect 11920 24731 11932 26307
rect 11874 24719 11932 24731
rect 12002 26307 12060 26319
rect 12002 24731 12014 26307
rect 12048 24731 12060 26307
rect 12002 24719 12060 24731
rect 12130 26307 12188 26319
rect 12130 24731 12142 26307
rect 12176 24731 12188 26307
rect 12130 24719 12188 24731
rect 12258 26307 12316 26319
rect 12258 24731 12270 26307
rect 12304 24731 12316 26307
rect 12258 24719 12316 24731
rect 19568 24707 19626 24719
rect 19568 23131 19580 24707
rect 19614 23131 19626 24707
rect 19568 23119 19626 23131
rect 19696 24707 19754 24719
rect 19696 23131 19708 24707
rect 19742 23131 19754 24707
rect 19696 23119 19754 23131
rect 19824 24707 19882 24719
rect 19824 23131 19836 24707
rect 19870 23131 19882 24707
rect 19824 23119 19882 23131
rect 19952 24707 20010 24719
rect 19952 23131 19964 24707
rect 19998 23131 20010 24707
rect 19952 23119 20010 23131
rect 20080 24707 20138 24719
rect 20080 23131 20092 24707
rect 20126 23131 20138 24707
rect 20080 23119 20138 23131
rect 20208 24707 20266 24719
rect 20208 23131 20220 24707
rect 20254 23131 20266 24707
rect 20208 23119 20266 23131
rect 20808 26307 20866 26319
rect 20808 24731 20820 26307
rect 20854 24731 20866 26307
rect 20808 24719 20866 24731
rect 20936 26307 20994 26319
rect 20936 24731 20948 26307
rect 20982 24731 20994 26307
rect 20936 24719 20994 24731
rect 21064 26307 21122 26319
rect 21064 24731 21076 26307
rect 21110 24731 21122 26307
rect 21064 24719 21122 24731
rect 21192 26307 21250 26319
rect 21192 24731 21204 26307
rect 21238 24731 21250 26307
rect 21192 24719 21250 24731
rect 21320 26307 21378 26319
rect 21320 24731 21332 26307
rect 21366 24731 21378 26307
rect 21320 24719 21378 24731
rect 21448 26307 21506 26319
rect 21448 24731 21460 26307
rect 21494 24731 21506 26307
rect 21448 24719 21506 24731
<< mvndiff >>
rect 31425 25775 33425 25787
rect 31425 25741 31437 25775
rect 33413 25741 33425 25775
rect 31425 25729 33425 25741
rect 31425 25617 33425 25629
rect 31425 25583 31437 25617
rect 33413 25583 33425 25617
rect 31425 25571 33425 25583
rect 30342 20238 30400 20250
rect 30342 19662 30354 20238
rect 30388 19662 30400 20238
rect 30342 19650 30400 19662
rect 30600 20238 30658 20250
rect 30600 19662 30612 20238
rect 30646 19662 30658 20238
rect 30600 19650 30658 19662
rect 30858 20238 30916 20250
rect 30858 19662 30870 20238
rect 30904 19662 30916 20238
rect 30858 19650 30916 19662
rect 31116 20238 31174 20250
rect 31116 19662 31128 20238
rect 31162 19662 31174 20238
rect 31116 19650 31174 19662
rect 31374 20238 31432 20250
rect 31374 19662 31386 20238
rect 31420 19662 31432 20238
rect 31374 19650 31432 19662
rect 31632 20238 31690 20250
rect 31632 19662 31644 20238
rect 31678 19662 31690 20238
rect 31632 19650 31690 19662
rect 31890 20238 31948 20250
rect 31890 19662 31902 20238
rect 31936 19662 31948 20238
rect 31890 19650 31948 19662
rect 32148 20238 32206 20250
rect 32148 19662 32160 20238
rect 32194 19662 32206 20238
rect 32148 19650 32206 19662
rect 33472 19438 33530 19450
rect 33472 18062 33484 19438
rect 33518 18062 33530 19438
rect 33472 18050 33530 18062
rect 33630 19438 33688 19450
rect 33630 18062 33642 19438
rect 33676 18062 33688 19438
rect 33630 18050 33688 18062
rect 33472 17538 33530 17550
rect 33472 16162 33484 17538
rect 33518 16162 33530 17538
rect 33472 16150 33530 16162
rect 33630 17538 33688 17550
rect 33630 16162 33642 17538
rect 33676 16162 33688 17538
rect 33630 16150 33688 16162
<< mvpdiff >>
rect 28760 19025 28818 19037
rect 28760 18449 28772 19025
rect 28806 18449 28818 19025
rect 28760 18437 28818 18449
rect 29018 19025 29076 19037
rect 29018 18449 29030 19025
rect 29064 18449 29076 19025
rect 29018 18437 29076 18449
rect 29276 19025 29334 19037
rect 29276 18449 29288 19025
rect 29322 18449 29334 19025
rect 29276 18437 29334 18449
rect 29534 19025 29592 19037
rect 29534 18449 29546 19025
rect 29580 18449 29592 19025
rect 29534 18437 29592 18449
rect 29792 19025 29850 19037
rect 29792 18449 29804 19025
rect 29838 18449 29850 19025
rect 29792 18437 29850 18449
rect 30050 19025 30108 19037
rect 30050 18449 30062 19025
rect 30096 18449 30108 19025
rect 30050 18437 30108 18449
rect 30308 19025 30366 19037
rect 30308 18449 30320 19025
rect 30354 18449 30366 19025
rect 30308 18437 30366 18449
rect 30566 19025 30624 19037
rect 30566 18449 30578 19025
rect 30612 18449 30624 19025
rect 30566 18437 30624 18449
rect 30824 19025 30882 19037
rect 30824 18449 30836 19025
rect 30870 18449 30882 19025
rect 30824 18437 30882 18449
rect 31082 19025 31140 19037
rect 31082 18449 31094 19025
rect 31128 18449 31140 19025
rect 31082 18437 31140 18449
rect 31340 19025 31398 19037
rect 31340 18449 31352 19025
rect 31386 18449 31398 19025
rect 31340 18437 31398 18449
rect 31598 19025 31656 19037
rect 31598 18449 31610 19025
rect 31644 18449 31656 19025
rect 31598 18437 31656 18449
rect 31856 19025 31914 19037
rect 31856 18449 31868 19025
rect 31902 18449 31914 19025
rect 31856 18437 31914 18449
rect 32114 19025 32172 19037
rect 32114 18449 32126 19025
rect 32160 18449 32172 19025
rect 32114 18437 32172 18449
rect 30050 17905 30108 17917
rect 30050 17329 30062 17905
rect 30096 17329 30108 17905
rect 30050 17317 30108 17329
rect 30308 17905 30366 17917
rect 30308 17329 30320 17905
rect 30354 17329 30366 17905
rect 30308 17317 30366 17329
rect 30566 17905 30624 17917
rect 30566 17329 30578 17905
rect 30612 17329 30624 17905
rect 30566 17317 30624 17329
rect 30824 17905 30882 17917
rect 30824 17329 30836 17905
rect 30870 17329 30882 17905
rect 30824 17317 30882 17329
rect 31082 17905 31140 17917
rect 31082 17329 31094 17905
rect 31128 17329 31140 17905
rect 31082 17317 31140 17329
rect 31340 17905 31398 17917
rect 31340 17329 31352 17905
rect 31386 17329 31398 17905
rect 31340 17317 31398 17329
rect 31598 17905 31656 17917
rect 31598 17329 31610 17905
rect 31644 17329 31656 17905
rect 31598 17317 31656 17329
rect 31856 17905 31914 17917
rect 31856 17329 31868 17905
rect 31902 17329 31914 17905
rect 31856 17317 31914 17329
rect 32114 17905 32172 17917
rect 32114 17329 32126 17905
rect 32160 17329 32172 17905
rect 32114 17317 32172 17329
rect 32830 18445 32888 18457
rect 32830 18069 32842 18445
rect 32876 18069 32888 18445
rect 32830 18057 32888 18069
rect 32988 18445 33046 18457
rect 32988 18069 33000 18445
rect 33034 18069 33046 18445
rect 32988 18057 33046 18069
rect 30050 16775 30108 16787
rect 30050 16199 30062 16775
rect 30096 16199 30108 16775
rect 30050 16187 30108 16199
rect 30308 16775 30366 16787
rect 30308 16199 30320 16775
rect 30354 16199 30366 16775
rect 30308 16187 30366 16199
rect 30566 16775 30624 16787
rect 30566 16199 30578 16775
rect 30612 16199 30624 16775
rect 30566 16187 30624 16199
rect 30824 16775 30882 16787
rect 30824 16199 30836 16775
rect 30870 16199 30882 16775
rect 30824 16187 30882 16199
rect 31082 16775 31140 16787
rect 31082 16199 31094 16775
rect 31128 16199 31140 16775
rect 31082 16187 31140 16199
rect 31340 16775 31398 16787
rect 31340 16199 31352 16775
rect 31386 16199 31398 16775
rect 31340 16187 31398 16199
rect 31598 16775 31656 16787
rect 31598 16199 31610 16775
rect 31644 16199 31656 16775
rect 31598 16187 31656 16199
rect 31856 16775 31914 16787
rect 31856 16199 31868 16775
rect 31902 16199 31914 16775
rect 31856 16187 31914 16199
rect 32114 16775 32172 16787
rect 32114 16199 32126 16775
rect 32160 16199 32172 16775
rect 32114 16187 32172 16199
rect 32830 17525 32888 17537
rect 32830 17149 32842 17525
rect 32876 17149 32888 17525
rect 32830 17137 32888 17149
rect 32988 17525 33046 17537
rect 32988 17149 33000 17525
rect 33034 17149 33046 17525
rect 32988 17137 33046 17149
<< pdiffc >>
rect 1250 23131 1284 24707
rect 1378 23131 1412 24707
rect 1506 23131 1540 24707
rect 1634 23131 1668 24707
rect 1762 23131 1796 24707
rect 1890 23131 1924 24707
rect 2490 24731 2524 26307
rect 2618 24731 2652 26307
rect 2746 24731 2780 26307
rect 2874 24731 2908 26307
rect 3002 24731 3036 26307
rect 3130 24731 3164 26307
rect 10390 23131 10424 24707
rect 10518 23131 10552 24707
rect 10646 23131 10680 24707
rect 10774 23131 10808 24707
rect 10902 23131 10936 24707
rect 11030 23131 11064 24707
rect 11630 24731 11664 26307
rect 11758 24731 11792 26307
rect 11886 24731 11920 26307
rect 12014 24731 12048 26307
rect 12142 24731 12176 26307
rect 12270 24731 12304 26307
rect 19580 23131 19614 24707
rect 19708 23131 19742 24707
rect 19836 23131 19870 24707
rect 19964 23131 19998 24707
rect 20092 23131 20126 24707
rect 20220 23131 20254 24707
rect 20820 24731 20854 26307
rect 20948 24731 20982 26307
rect 21076 24731 21110 26307
rect 21204 24731 21238 26307
rect 21332 24731 21366 26307
rect 21460 24731 21494 26307
<< mvndiffc >>
rect 31437 25741 33413 25775
rect 31437 25583 33413 25617
rect 30354 19662 30388 20238
rect 30612 19662 30646 20238
rect 30870 19662 30904 20238
rect 31128 19662 31162 20238
rect 31386 19662 31420 20238
rect 31644 19662 31678 20238
rect 31902 19662 31936 20238
rect 32160 19662 32194 20238
rect 33484 18062 33518 19438
rect 33642 18062 33676 19438
rect 33484 16162 33518 17538
rect 33642 16162 33676 17538
<< mvpdiffc >>
rect 28772 18449 28806 19025
rect 29030 18449 29064 19025
rect 29288 18449 29322 19025
rect 29546 18449 29580 19025
rect 29804 18449 29838 19025
rect 30062 18449 30096 19025
rect 30320 18449 30354 19025
rect 30578 18449 30612 19025
rect 30836 18449 30870 19025
rect 31094 18449 31128 19025
rect 31352 18449 31386 19025
rect 31610 18449 31644 19025
rect 31868 18449 31902 19025
rect 32126 18449 32160 19025
rect 30062 17329 30096 17905
rect 30320 17329 30354 17905
rect 30578 17329 30612 17905
rect 30836 17329 30870 17905
rect 31094 17329 31128 17905
rect 31352 17329 31386 17905
rect 31610 17329 31644 17905
rect 31868 17329 31902 17905
rect 32126 17329 32160 17905
rect 32842 18069 32876 18445
rect 33000 18069 33034 18445
rect 30062 16199 30096 16775
rect 30320 16199 30354 16775
rect 30578 16199 30612 16775
rect 30836 16199 30870 16775
rect 31094 16199 31128 16775
rect 31352 16199 31386 16775
rect 31610 16199 31644 16775
rect 31868 16199 31902 16775
rect 32126 16199 32160 16775
rect 32842 17149 32876 17525
rect 33000 17149 33034 17525
<< nsubdiff >>
rect 2376 26468 2472 26502
rect 3182 26468 3278 26502
rect 2376 26406 2410 26468
rect 1136 24868 1232 24902
rect 1942 24868 2038 24902
rect 1136 24806 1170 24868
rect 2004 24806 2038 24868
rect 1136 22970 1170 23032
rect 3244 26406 3278 26468
rect 2376 24570 2410 24632
rect 11516 26468 11612 26502
rect 12322 26468 12418 26502
rect 11516 26406 11550 26468
rect 3244 24570 3278 24632
rect 2376 24536 2472 24570
rect 3182 24536 3278 24570
rect 10276 24868 10372 24902
rect 11082 24868 11178 24902
rect 10276 24806 10310 24868
rect 2004 22970 2038 23032
rect 1136 22936 1232 22970
rect 1942 22936 2038 22970
rect 11144 24806 11178 24868
rect 10276 22970 10310 23032
rect 12384 26406 12418 26468
rect 11516 24570 11550 24632
rect 20706 26468 20802 26502
rect 21512 26468 21608 26502
rect 20706 26406 20740 26468
rect 12384 24570 12418 24632
rect 11516 24536 11612 24570
rect 12322 24536 12418 24570
rect 19466 24868 19562 24902
rect 20272 24868 20368 24902
rect 19466 24806 19500 24868
rect 11144 22970 11178 23032
rect 10276 22936 10372 22970
rect 11082 22936 11178 22970
rect 20334 24806 20368 24868
rect 19466 22970 19500 23032
rect 21574 26406 21608 26468
rect 20706 24570 20740 24632
rect 21574 24570 21608 24632
rect 20706 24536 20802 24570
rect 21512 24536 21608 24570
rect 20334 22970 20368 23032
rect 19466 22936 19562 22970
rect 20272 22936 20368 22970
<< mvpsubdiff >>
rect 31203 25909 33647 25921
rect 31203 25875 31311 25909
rect 33539 25875 33647 25909
rect 31203 25863 33647 25875
rect 31203 25813 31261 25863
rect 31203 25545 31215 25813
rect 31249 25545 31261 25813
rect 33589 25813 33647 25863
rect 31203 25495 31261 25545
rect 33589 25545 33601 25813
rect 33635 25545 33647 25813
rect 33589 25495 33647 25545
rect 31203 25483 33647 25495
rect 31203 25449 31311 25483
rect 33539 25449 33647 25483
rect 31203 25437 33647 25449
rect 30208 20460 32340 20472
rect 30208 20426 30316 20460
rect 32232 20426 32340 20460
rect 30208 20414 32340 20426
rect 30208 20364 30266 20414
rect 30208 19536 30220 20364
rect 30254 19536 30266 20364
rect 32282 20364 32340 20414
rect 30208 19486 30266 19536
rect 32282 19536 32294 20364
rect 32328 19536 32340 20364
rect 32282 19486 32340 19536
rect 30208 19474 32340 19486
rect 30208 19440 30316 19474
rect 32232 19440 32340 19474
rect 30208 19428 32340 19440
rect 33338 19660 33822 19672
rect 33338 19626 33446 19660
rect 33714 19626 33822 19660
rect 33338 19614 33822 19626
rect 33338 19564 33396 19614
rect 33338 17936 33350 19564
rect 33384 17936 33396 19564
rect 33764 19564 33822 19614
rect 33338 17886 33396 17936
rect 33764 17936 33776 19564
rect 33810 17936 33822 19564
rect 33764 17886 33822 17936
rect 33338 17874 33822 17886
rect 33338 17840 33446 17874
rect 33714 17840 33822 17874
rect 33338 17828 33822 17840
rect 33338 17760 33822 17772
rect 33338 17726 33446 17760
rect 33714 17726 33822 17760
rect 33338 17714 33822 17726
rect 33338 17664 33396 17714
rect 33338 16036 33350 17664
rect 33384 16036 33396 17664
rect 33764 17664 33822 17714
rect 33338 15986 33396 16036
rect 33764 16036 33776 17664
rect 33810 16036 33822 17664
rect 33764 15986 33822 16036
rect 33338 15974 33822 15986
rect 33338 15940 33446 15974
rect 33714 15940 33822 15974
rect 33338 15928 33822 15940
<< mvnsubdiff >>
rect 28626 19256 32306 19268
rect 28626 19222 28734 19256
rect 32198 19222 32306 19256
rect 28626 19210 32306 19222
rect 28626 19160 28684 19210
rect 28626 18314 28638 19160
rect 28672 18314 28684 19160
rect 32248 19160 32306 19210
rect 28626 18264 28684 18314
rect 32248 18314 32260 19160
rect 32294 18314 32306 19160
rect 32248 18264 32306 18314
rect 28626 18252 32306 18264
rect 28626 18218 28734 18252
rect 32198 18218 32306 18252
rect 28626 18206 32306 18218
rect 32696 18676 33180 18688
rect 32696 18642 32804 18676
rect 33072 18642 33180 18676
rect 32696 18630 33180 18642
rect 32696 18580 32754 18630
rect 29916 18136 32306 18148
rect 29916 18102 30024 18136
rect 32198 18102 32306 18136
rect 29916 18090 32306 18102
rect 29916 18040 29974 18090
rect 29916 17194 29928 18040
rect 29962 17194 29974 18040
rect 32248 18040 32306 18090
rect 29916 17144 29974 17194
rect 32248 17194 32260 18040
rect 32294 17194 32306 18040
rect 32696 17934 32708 18580
rect 32742 17934 32754 18580
rect 33122 18580 33180 18630
rect 32696 17884 32754 17934
rect 33122 17934 33134 18580
rect 33168 17934 33180 18580
rect 33122 17884 33180 17934
rect 32696 17872 33180 17884
rect 32696 17838 32804 17872
rect 33072 17838 33180 17872
rect 32696 17826 33180 17838
rect 32248 17144 32306 17194
rect 29916 17132 32306 17144
rect 29916 17098 30024 17132
rect 32198 17098 32306 17132
rect 29916 17086 32306 17098
rect 32696 17756 33180 17768
rect 32696 17722 32804 17756
rect 33072 17722 33180 17756
rect 32696 17710 33180 17722
rect 32696 17660 32754 17710
rect 29916 17006 32306 17018
rect 29916 16972 30024 17006
rect 32198 16972 32306 17006
rect 29916 16960 32306 16972
rect 29916 16910 29974 16960
rect 29916 16064 29928 16910
rect 29962 16064 29974 16910
rect 32248 16910 32306 16960
rect 29916 16014 29974 16064
rect 32248 16064 32260 16910
rect 32294 16064 32306 16910
rect 32696 17014 32708 17660
rect 32742 17014 32754 17660
rect 33122 17660 33180 17710
rect 32696 16964 32754 17014
rect 33122 17014 33134 17660
rect 33168 17014 33180 17660
rect 33122 16964 33180 17014
rect 32696 16952 33180 16964
rect 32696 16918 32804 16952
rect 33072 16918 33180 16952
rect 32696 16906 33180 16918
rect 32248 16014 32306 16064
rect 29916 16002 32306 16014
rect 29916 15968 30024 16002
rect 32198 15968 32306 16002
rect 29916 15956 32306 15968
<< nsubdiffcont >>
rect 2472 26468 3182 26502
rect 1232 24868 1942 24902
rect 1136 23032 1170 24806
rect 2004 23032 2038 24806
rect 2376 24632 2410 26406
rect 3244 24632 3278 26406
rect 11612 26468 12322 26502
rect 2472 24536 3182 24570
rect 10372 24868 11082 24902
rect 1232 22936 1942 22970
rect 10276 23032 10310 24806
rect 11144 23032 11178 24806
rect 11516 24632 11550 26406
rect 12384 24632 12418 26406
rect 20802 26468 21512 26502
rect 11612 24536 12322 24570
rect 19562 24868 20272 24902
rect 10372 22936 11082 22970
rect 19466 23032 19500 24806
rect 20334 23032 20368 24806
rect 20706 24632 20740 26406
rect 21574 24632 21608 26406
rect 20802 24536 21512 24570
rect 19562 22936 20272 22970
<< mvpsubdiffcont >>
rect 31311 25875 33539 25909
rect 31215 25545 31249 25813
rect 33601 25545 33635 25813
rect 31311 25449 33539 25483
rect 30316 20426 32232 20460
rect 30220 19536 30254 20364
rect 32294 19536 32328 20364
rect 30316 19440 32232 19474
rect 33446 19626 33714 19660
rect 33350 17936 33384 19564
rect 33776 17936 33810 19564
rect 33446 17840 33714 17874
rect 33446 17726 33714 17760
rect 33350 16036 33384 17664
rect 33776 16036 33810 17664
rect 33446 15940 33714 15974
<< mvnsubdiffcont >>
rect 28734 19222 32198 19256
rect 28638 18314 28672 19160
rect 32260 18314 32294 19160
rect 28734 18218 32198 18252
rect 32804 18642 33072 18676
rect 30024 18102 32198 18136
rect 29928 17194 29962 18040
rect 32260 17194 32294 18040
rect 32708 17934 32742 18580
rect 33134 17934 33168 18580
rect 32804 17838 33072 17872
rect 30024 17098 32198 17132
rect 32804 17722 33072 17756
rect 30024 16972 32198 17006
rect 29928 16064 29962 16910
rect 32260 16064 32294 16910
rect 32708 17014 32742 17660
rect 33134 17014 33168 17660
rect 32804 16918 33072 16952
rect 30024 15968 32198 16002
<< poly >>
rect 1296 24800 1366 24816
rect 1296 24766 1312 24800
rect 1350 24766 1366 24800
rect 1296 24719 1366 24766
rect 1424 24800 1494 24816
rect 1424 24766 1440 24800
rect 1478 24766 1494 24800
rect 1424 24719 1494 24766
rect 1552 24800 1622 24816
rect 1552 24766 1568 24800
rect 1606 24766 1622 24800
rect 1552 24719 1622 24766
rect 1680 24800 1750 24816
rect 1680 24766 1696 24800
rect 1734 24766 1750 24800
rect 1680 24719 1750 24766
rect 1808 24800 1878 24816
rect 1808 24766 1824 24800
rect 1862 24766 1878 24800
rect 1808 24719 1878 24766
rect 1296 23072 1366 23119
rect 1296 23038 1312 23072
rect 1350 23038 1366 23072
rect 1296 23022 1366 23038
rect 1424 23072 1494 23119
rect 1424 23038 1440 23072
rect 1478 23038 1494 23072
rect 1424 23022 1494 23038
rect 1552 23072 1622 23119
rect 1552 23038 1568 23072
rect 1606 23038 1622 23072
rect 1552 23022 1622 23038
rect 1680 23072 1750 23119
rect 1680 23038 1696 23072
rect 1734 23038 1750 23072
rect 1680 23022 1750 23038
rect 1808 23072 1878 23119
rect 1808 23038 1824 23072
rect 1862 23038 1878 23072
rect 1808 23022 1878 23038
rect 2536 26400 2606 26416
rect 2536 26366 2552 26400
rect 2590 26366 2606 26400
rect 2536 26319 2606 26366
rect 2664 26400 2734 26416
rect 2664 26366 2680 26400
rect 2718 26366 2734 26400
rect 2664 26319 2734 26366
rect 2792 26400 2862 26416
rect 2792 26366 2808 26400
rect 2846 26366 2862 26400
rect 2792 26319 2862 26366
rect 2920 26400 2990 26416
rect 2920 26366 2936 26400
rect 2974 26366 2990 26400
rect 2920 26319 2990 26366
rect 3048 26400 3118 26416
rect 3048 26366 3064 26400
rect 3102 26366 3118 26400
rect 3048 26319 3118 26366
rect 2536 24672 2606 24719
rect 2536 24638 2552 24672
rect 2590 24638 2606 24672
rect 2536 24622 2606 24638
rect 2664 24672 2734 24719
rect 2664 24638 2680 24672
rect 2718 24638 2734 24672
rect 2664 24622 2734 24638
rect 2792 24672 2862 24719
rect 2792 24638 2808 24672
rect 2846 24638 2862 24672
rect 2792 24622 2862 24638
rect 2920 24672 2990 24719
rect 2920 24638 2936 24672
rect 2974 24638 2990 24672
rect 2920 24622 2990 24638
rect 3048 24672 3118 24719
rect 3048 24638 3064 24672
rect 3102 24638 3118 24672
rect 3048 24622 3118 24638
rect 10436 24800 10506 24816
rect 10436 24766 10452 24800
rect 10490 24766 10506 24800
rect 10436 24719 10506 24766
rect 10564 24800 10634 24816
rect 10564 24766 10580 24800
rect 10618 24766 10634 24800
rect 10564 24719 10634 24766
rect 10692 24800 10762 24816
rect 10692 24766 10708 24800
rect 10746 24766 10762 24800
rect 10692 24719 10762 24766
rect 10820 24800 10890 24816
rect 10820 24766 10836 24800
rect 10874 24766 10890 24800
rect 10820 24719 10890 24766
rect 10948 24800 11018 24816
rect 10948 24766 10964 24800
rect 11002 24766 11018 24800
rect 10948 24719 11018 24766
rect 10436 23072 10506 23119
rect 10436 23038 10452 23072
rect 10490 23038 10506 23072
rect 10436 23022 10506 23038
rect 10564 23072 10634 23119
rect 10564 23038 10580 23072
rect 10618 23038 10634 23072
rect 10564 23022 10634 23038
rect 10692 23072 10762 23119
rect 10692 23038 10708 23072
rect 10746 23038 10762 23072
rect 10692 23022 10762 23038
rect 10820 23072 10890 23119
rect 10820 23038 10836 23072
rect 10874 23038 10890 23072
rect 10820 23022 10890 23038
rect 10948 23072 11018 23119
rect 10948 23038 10964 23072
rect 11002 23038 11018 23072
rect 10948 23022 11018 23038
rect 11676 26400 11746 26416
rect 11676 26366 11692 26400
rect 11730 26366 11746 26400
rect 11676 26319 11746 26366
rect 11804 26400 11874 26416
rect 11804 26366 11820 26400
rect 11858 26366 11874 26400
rect 11804 26319 11874 26366
rect 11932 26400 12002 26416
rect 11932 26366 11948 26400
rect 11986 26366 12002 26400
rect 11932 26319 12002 26366
rect 12060 26400 12130 26416
rect 12060 26366 12076 26400
rect 12114 26366 12130 26400
rect 12060 26319 12130 26366
rect 12188 26400 12258 26416
rect 12188 26366 12204 26400
rect 12242 26366 12258 26400
rect 12188 26319 12258 26366
rect 11676 24672 11746 24719
rect 11676 24638 11692 24672
rect 11730 24638 11746 24672
rect 11676 24622 11746 24638
rect 11804 24672 11874 24719
rect 11804 24638 11820 24672
rect 11858 24638 11874 24672
rect 11804 24622 11874 24638
rect 11932 24672 12002 24719
rect 11932 24638 11948 24672
rect 11986 24638 12002 24672
rect 11932 24622 12002 24638
rect 12060 24672 12130 24719
rect 12060 24638 12076 24672
rect 12114 24638 12130 24672
rect 12060 24622 12130 24638
rect 12188 24672 12258 24719
rect 12188 24638 12204 24672
rect 12242 24638 12258 24672
rect 12188 24622 12258 24638
rect 19626 24800 19696 24816
rect 19626 24766 19642 24800
rect 19680 24766 19696 24800
rect 19626 24719 19696 24766
rect 19754 24800 19824 24816
rect 19754 24766 19770 24800
rect 19808 24766 19824 24800
rect 19754 24719 19824 24766
rect 19882 24800 19952 24816
rect 19882 24766 19898 24800
rect 19936 24766 19952 24800
rect 19882 24719 19952 24766
rect 20010 24800 20080 24816
rect 20010 24766 20026 24800
rect 20064 24766 20080 24800
rect 20010 24719 20080 24766
rect 20138 24800 20208 24816
rect 20138 24766 20154 24800
rect 20192 24766 20208 24800
rect 20138 24719 20208 24766
rect 19626 23072 19696 23119
rect 19626 23038 19642 23072
rect 19680 23038 19696 23072
rect 19626 23022 19696 23038
rect 19754 23072 19824 23119
rect 19754 23038 19770 23072
rect 19808 23038 19824 23072
rect 19754 23022 19824 23038
rect 19882 23072 19952 23119
rect 19882 23038 19898 23072
rect 19936 23038 19952 23072
rect 19882 23022 19952 23038
rect 20010 23072 20080 23119
rect 20010 23038 20026 23072
rect 20064 23038 20080 23072
rect 20010 23022 20080 23038
rect 20138 23072 20208 23119
rect 20138 23038 20154 23072
rect 20192 23038 20208 23072
rect 20138 23022 20208 23038
rect 20866 26400 20936 26416
rect 20866 26366 20882 26400
rect 20920 26366 20936 26400
rect 20866 26319 20936 26366
rect 20994 26400 21064 26416
rect 20994 26366 21010 26400
rect 21048 26366 21064 26400
rect 20994 26319 21064 26366
rect 21122 26400 21192 26416
rect 21122 26366 21138 26400
rect 21176 26366 21192 26400
rect 21122 26319 21192 26366
rect 21250 26400 21320 26416
rect 21250 26366 21266 26400
rect 21304 26366 21320 26400
rect 21250 26319 21320 26366
rect 21378 26400 21448 26416
rect 21378 26366 21394 26400
rect 21432 26366 21448 26400
rect 21378 26319 21448 26366
rect 20866 24672 20936 24719
rect 20866 24638 20882 24672
rect 20920 24638 20936 24672
rect 20866 24622 20936 24638
rect 20994 24672 21064 24719
rect 20994 24638 21010 24672
rect 21048 24638 21064 24672
rect 20994 24622 21064 24638
rect 21122 24672 21192 24719
rect 21122 24638 21138 24672
rect 21176 24638 21192 24672
rect 21122 24622 21192 24638
rect 21250 24672 21320 24719
rect 21250 24638 21266 24672
rect 21304 24638 21320 24672
rect 21250 24622 21320 24638
rect 21378 24672 21448 24719
rect 21378 24638 21394 24672
rect 21432 24638 21448 24672
rect 21378 24622 21448 24638
rect 31337 25713 31425 25729
rect 31337 25645 31353 25713
rect 31387 25645 31425 25713
rect 31337 25629 31425 25645
rect 33425 25713 33513 25729
rect 33425 25645 33463 25713
rect 33497 25645 33513 25713
rect 33425 25629 33513 25645
rect 30400 20322 30600 20338
rect 30400 20288 30416 20322
rect 30584 20288 30600 20322
rect 30400 20250 30600 20288
rect 30658 20322 30858 20338
rect 30658 20288 30674 20322
rect 30842 20288 30858 20322
rect 30658 20250 30858 20288
rect 30916 20322 31116 20338
rect 30916 20288 30932 20322
rect 31100 20288 31116 20322
rect 30916 20250 31116 20288
rect 31174 20322 31374 20338
rect 31174 20288 31190 20322
rect 31358 20288 31374 20322
rect 31174 20250 31374 20288
rect 31432 20322 31632 20338
rect 31432 20288 31448 20322
rect 31616 20288 31632 20322
rect 31432 20250 31632 20288
rect 31690 20322 31890 20338
rect 31690 20288 31706 20322
rect 31874 20288 31890 20322
rect 31690 20250 31890 20288
rect 31948 20322 32148 20338
rect 31948 20288 31964 20322
rect 32132 20288 32148 20322
rect 31948 20250 32148 20288
rect 30400 19612 30600 19650
rect 30400 19578 30416 19612
rect 30584 19578 30600 19612
rect 30400 19562 30600 19578
rect 30658 19612 30858 19650
rect 30658 19578 30674 19612
rect 30842 19578 30858 19612
rect 30658 19562 30858 19578
rect 30916 19612 31116 19650
rect 30916 19578 30932 19612
rect 31100 19578 31116 19612
rect 30916 19562 31116 19578
rect 31174 19612 31374 19650
rect 31174 19578 31190 19612
rect 31358 19578 31374 19612
rect 31174 19562 31374 19578
rect 31432 19612 31632 19650
rect 31432 19578 31448 19612
rect 31616 19578 31632 19612
rect 31432 19562 31632 19578
rect 31690 19612 31890 19650
rect 31690 19578 31706 19612
rect 31874 19578 31890 19612
rect 31690 19562 31890 19578
rect 31948 19612 32148 19650
rect 31948 19578 31964 19612
rect 32132 19578 32148 19612
rect 31948 19562 32148 19578
rect 28818 19118 29018 19134
rect 28818 19084 28834 19118
rect 29002 19084 29018 19118
rect 28818 19037 29018 19084
rect 29076 19118 29276 19134
rect 29076 19084 29092 19118
rect 29260 19084 29276 19118
rect 29076 19037 29276 19084
rect 29334 19118 29534 19134
rect 29334 19084 29350 19118
rect 29518 19084 29534 19118
rect 29334 19037 29534 19084
rect 29592 19118 29792 19134
rect 29592 19084 29608 19118
rect 29776 19084 29792 19118
rect 29592 19037 29792 19084
rect 29850 19118 30050 19134
rect 29850 19084 29866 19118
rect 30034 19084 30050 19118
rect 29850 19037 30050 19084
rect 30108 19118 30308 19134
rect 30108 19084 30124 19118
rect 30292 19084 30308 19118
rect 30108 19037 30308 19084
rect 30366 19118 30566 19134
rect 30366 19084 30382 19118
rect 30550 19084 30566 19118
rect 30366 19037 30566 19084
rect 30624 19118 30824 19134
rect 30624 19084 30640 19118
rect 30808 19084 30824 19118
rect 30624 19037 30824 19084
rect 30882 19118 31082 19134
rect 30882 19084 30898 19118
rect 31066 19084 31082 19118
rect 30882 19037 31082 19084
rect 31140 19118 31340 19134
rect 31140 19084 31156 19118
rect 31324 19084 31340 19118
rect 31140 19037 31340 19084
rect 31398 19118 31598 19134
rect 31398 19084 31414 19118
rect 31582 19084 31598 19118
rect 31398 19037 31598 19084
rect 31656 19118 31856 19134
rect 31656 19084 31672 19118
rect 31840 19084 31856 19118
rect 31656 19037 31856 19084
rect 31914 19118 32114 19134
rect 31914 19084 31930 19118
rect 32098 19084 32114 19118
rect 31914 19037 32114 19084
rect 28818 18390 29018 18437
rect 28818 18356 28834 18390
rect 29002 18356 29018 18390
rect 28818 18340 29018 18356
rect 29076 18390 29276 18437
rect 29076 18356 29092 18390
rect 29260 18356 29276 18390
rect 29076 18340 29276 18356
rect 29334 18390 29534 18437
rect 29334 18356 29350 18390
rect 29518 18356 29534 18390
rect 29334 18340 29534 18356
rect 29592 18390 29792 18437
rect 29592 18356 29608 18390
rect 29776 18356 29792 18390
rect 29592 18340 29792 18356
rect 29850 18390 30050 18437
rect 29850 18356 29866 18390
rect 30034 18356 30050 18390
rect 29850 18340 30050 18356
rect 30108 18390 30308 18437
rect 30108 18356 30124 18390
rect 30292 18356 30308 18390
rect 30108 18340 30308 18356
rect 30366 18390 30566 18437
rect 30366 18356 30382 18390
rect 30550 18356 30566 18390
rect 30366 18340 30566 18356
rect 30624 18390 30824 18437
rect 30624 18356 30640 18390
rect 30808 18356 30824 18390
rect 30624 18340 30824 18356
rect 30882 18390 31082 18437
rect 30882 18356 30898 18390
rect 31066 18356 31082 18390
rect 30882 18340 31082 18356
rect 31140 18390 31340 18437
rect 31140 18356 31156 18390
rect 31324 18356 31340 18390
rect 31140 18340 31340 18356
rect 31398 18390 31598 18437
rect 31398 18356 31414 18390
rect 31582 18356 31598 18390
rect 31398 18340 31598 18356
rect 31656 18390 31856 18437
rect 31656 18356 31672 18390
rect 31840 18356 31856 18390
rect 31656 18340 31856 18356
rect 31914 18390 32114 18437
rect 31914 18356 31930 18390
rect 32098 18356 32114 18390
rect 31914 18340 32114 18356
rect 30108 17998 30308 18014
rect 30108 17964 30124 17998
rect 30292 17964 30308 17998
rect 30108 17917 30308 17964
rect 30366 17998 30566 18014
rect 30366 17964 30382 17998
rect 30550 17964 30566 17998
rect 30366 17917 30566 17964
rect 30624 17998 30824 18014
rect 30624 17964 30640 17998
rect 30808 17964 30824 17998
rect 30624 17917 30824 17964
rect 30882 17998 31082 18014
rect 30882 17964 30898 17998
rect 31066 17964 31082 17998
rect 30882 17917 31082 17964
rect 31140 17998 31340 18014
rect 31140 17964 31156 17998
rect 31324 17964 31340 17998
rect 31140 17917 31340 17964
rect 31398 17998 31598 18014
rect 31398 17964 31414 17998
rect 31582 17964 31598 17998
rect 31398 17917 31598 17964
rect 31656 17998 31856 18014
rect 31656 17964 31672 17998
rect 31840 17964 31856 17998
rect 31656 17917 31856 17964
rect 31914 17998 32114 18014
rect 31914 17964 31930 17998
rect 32098 17964 32114 17998
rect 31914 17917 32114 17964
rect 30108 17270 30308 17317
rect 30108 17236 30124 17270
rect 30292 17236 30308 17270
rect 30108 17220 30308 17236
rect 30366 17270 30566 17317
rect 30366 17236 30382 17270
rect 30550 17236 30566 17270
rect 30366 17220 30566 17236
rect 30624 17270 30824 17317
rect 30624 17236 30640 17270
rect 30808 17236 30824 17270
rect 30624 17220 30824 17236
rect 30882 17270 31082 17317
rect 30882 17236 30898 17270
rect 31066 17236 31082 17270
rect 30882 17220 31082 17236
rect 31140 17270 31340 17317
rect 31140 17236 31156 17270
rect 31324 17236 31340 17270
rect 31140 17220 31340 17236
rect 31398 17270 31598 17317
rect 31398 17236 31414 17270
rect 31582 17236 31598 17270
rect 31398 17220 31598 17236
rect 31656 17270 31856 17317
rect 31656 17236 31672 17270
rect 31840 17236 31856 17270
rect 31656 17220 31856 17236
rect 31914 17270 32114 17317
rect 31914 17236 31930 17270
rect 32098 17236 32114 17270
rect 31914 17220 32114 17236
rect 32888 18538 32988 18554
rect 32888 18504 32904 18538
rect 32972 18504 32988 18538
rect 32888 18457 32988 18504
rect 32888 18010 32988 18057
rect 32888 17976 32904 18010
rect 32972 17976 32988 18010
rect 32888 17960 32988 17976
rect 33530 19522 33630 19538
rect 33530 19488 33546 19522
rect 33614 19488 33630 19522
rect 33530 19450 33630 19488
rect 33530 18012 33630 18050
rect 33530 17978 33546 18012
rect 33614 17978 33630 18012
rect 33530 17962 33630 17978
rect 30108 16868 30308 16884
rect 30108 16834 30124 16868
rect 30292 16834 30308 16868
rect 30108 16787 30308 16834
rect 30366 16868 30566 16884
rect 30366 16834 30382 16868
rect 30550 16834 30566 16868
rect 30366 16787 30566 16834
rect 30624 16868 30824 16884
rect 30624 16834 30640 16868
rect 30808 16834 30824 16868
rect 30624 16787 30824 16834
rect 30882 16868 31082 16884
rect 30882 16834 30898 16868
rect 31066 16834 31082 16868
rect 30882 16787 31082 16834
rect 31140 16868 31340 16884
rect 31140 16834 31156 16868
rect 31324 16834 31340 16868
rect 31140 16787 31340 16834
rect 31398 16868 31598 16884
rect 31398 16834 31414 16868
rect 31582 16834 31598 16868
rect 31398 16787 31598 16834
rect 31656 16868 31856 16884
rect 31656 16834 31672 16868
rect 31840 16834 31856 16868
rect 31656 16787 31856 16834
rect 31914 16868 32114 16884
rect 31914 16834 31930 16868
rect 32098 16834 32114 16868
rect 31914 16787 32114 16834
rect 30108 16140 30308 16187
rect 30108 16106 30124 16140
rect 30292 16106 30308 16140
rect 30108 16090 30308 16106
rect 30366 16140 30566 16187
rect 30366 16106 30382 16140
rect 30550 16106 30566 16140
rect 30366 16090 30566 16106
rect 30624 16140 30824 16187
rect 30624 16106 30640 16140
rect 30808 16106 30824 16140
rect 30624 16090 30824 16106
rect 30882 16140 31082 16187
rect 30882 16106 30898 16140
rect 31066 16106 31082 16140
rect 30882 16090 31082 16106
rect 31140 16140 31340 16187
rect 31140 16106 31156 16140
rect 31324 16106 31340 16140
rect 31140 16090 31340 16106
rect 31398 16140 31598 16187
rect 31398 16106 31414 16140
rect 31582 16106 31598 16140
rect 31398 16090 31598 16106
rect 31656 16140 31856 16187
rect 31656 16106 31672 16140
rect 31840 16106 31856 16140
rect 31656 16090 31856 16106
rect 31914 16140 32114 16187
rect 31914 16106 31930 16140
rect 32098 16106 32114 16140
rect 31914 16090 32114 16106
rect 32888 17618 32988 17634
rect 32888 17584 32904 17618
rect 32972 17584 32988 17618
rect 32888 17537 32988 17584
rect 32888 17090 32988 17137
rect 32888 17056 32904 17090
rect 32972 17056 32988 17090
rect 32888 17040 32988 17056
rect 33530 17622 33630 17638
rect 33530 17588 33546 17622
rect 33614 17588 33630 17622
rect 33530 17550 33630 17588
rect 33530 16112 33630 16150
rect 33530 16078 33546 16112
rect 33614 16078 33630 16112
rect 33530 16062 33630 16078
<< polycont >>
rect 1312 24766 1350 24800
rect 1440 24766 1478 24800
rect 1568 24766 1606 24800
rect 1696 24766 1734 24800
rect 1824 24766 1862 24800
rect 1312 23038 1350 23072
rect 1440 23038 1478 23072
rect 1568 23038 1606 23072
rect 1696 23038 1734 23072
rect 1824 23038 1862 23072
rect 2552 26366 2590 26400
rect 2680 26366 2718 26400
rect 2808 26366 2846 26400
rect 2936 26366 2974 26400
rect 3064 26366 3102 26400
rect 2552 24638 2590 24672
rect 2680 24638 2718 24672
rect 2808 24638 2846 24672
rect 2936 24638 2974 24672
rect 3064 24638 3102 24672
rect 10452 24766 10490 24800
rect 10580 24766 10618 24800
rect 10708 24766 10746 24800
rect 10836 24766 10874 24800
rect 10964 24766 11002 24800
rect 10452 23038 10490 23072
rect 10580 23038 10618 23072
rect 10708 23038 10746 23072
rect 10836 23038 10874 23072
rect 10964 23038 11002 23072
rect 11692 26366 11730 26400
rect 11820 26366 11858 26400
rect 11948 26366 11986 26400
rect 12076 26366 12114 26400
rect 12204 26366 12242 26400
rect 11692 24638 11730 24672
rect 11820 24638 11858 24672
rect 11948 24638 11986 24672
rect 12076 24638 12114 24672
rect 12204 24638 12242 24672
rect 19642 24766 19680 24800
rect 19770 24766 19808 24800
rect 19898 24766 19936 24800
rect 20026 24766 20064 24800
rect 20154 24766 20192 24800
rect 19642 23038 19680 23072
rect 19770 23038 19808 23072
rect 19898 23038 19936 23072
rect 20026 23038 20064 23072
rect 20154 23038 20192 23072
rect 20882 26366 20920 26400
rect 21010 26366 21048 26400
rect 21138 26366 21176 26400
rect 21266 26366 21304 26400
rect 21394 26366 21432 26400
rect 20882 24638 20920 24672
rect 21010 24638 21048 24672
rect 21138 24638 21176 24672
rect 21266 24638 21304 24672
rect 21394 24638 21432 24672
rect 31353 25645 31387 25713
rect 33463 25645 33497 25713
rect 30416 20288 30584 20322
rect 30674 20288 30842 20322
rect 30932 20288 31100 20322
rect 31190 20288 31358 20322
rect 31448 20288 31616 20322
rect 31706 20288 31874 20322
rect 31964 20288 32132 20322
rect 30416 19578 30584 19612
rect 30674 19578 30842 19612
rect 30932 19578 31100 19612
rect 31190 19578 31358 19612
rect 31448 19578 31616 19612
rect 31706 19578 31874 19612
rect 31964 19578 32132 19612
rect 28834 19084 29002 19118
rect 29092 19084 29260 19118
rect 29350 19084 29518 19118
rect 29608 19084 29776 19118
rect 29866 19084 30034 19118
rect 30124 19084 30292 19118
rect 30382 19084 30550 19118
rect 30640 19084 30808 19118
rect 30898 19084 31066 19118
rect 31156 19084 31324 19118
rect 31414 19084 31582 19118
rect 31672 19084 31840 19118
rect 31930 19084 32098 19118
rect 28834 18356 29002 18390
rect 29092 18356 29260 18390
rect 29350 18356 29518 18390
rect 29608 18356 29776 18390
rect 29866 18356 30034 18390
rect 30124 18356 30292 18390
rect 30382 18356 30550 18390
rect 30640 18356 30808 18390
rect 30898 18356 31066 18390
rect 31156 18356 31324 18390
rect 31414 18356 31582 18390
rect 31672 18356 31840 18390
rect 31930 18356 32098 18390
rect 30124 17964 30292 17998
rect 30382 17964 30550 17998
rect 30640 17964 30808 17998
rect 30898 17964 31066 17998
rect 31156 17964 31324 17998
rect 31414 17964 31582 17998
rect 31672 17964 31840 17998
rect 31930 17964 32098 17998
rect 30124 17236 30292 17270
rect 30382 17236 30550 17270
rect 30640 17236 30808 17270
rect 30898 17236 31066 17270
rect 31156 17236 31324 17270
rect 31414 17236 31582 17270
rect 31672 17236 31840 17270
rect 31930 17236 32098 17270
rect 32904 18504 32972 18538
rect 32904 17976 32972 18010
rect 33546 19488 33614 19522
rect 33546 17978 33614 18012
rect 30124 16834 30292 16868
rect 30382 16834 30550 16868
rect 30640 16834 30808 16868
rect 30898 16834 31066 16868
rect 31156 16834 31324 16868
rect 31414 16834 31582 16868
rect 31672 16834 31840 16868
rect 31930 16834 32098 16868
rect 30124 16106 30292 16140
rect 30382 16106 30550 16140
rect 30640 16106 30808 16140
rect 30898 16106 31066 16140
rect 31156 16106 31324 16140
rect 31414 16106 31582 16140
rect 31672 16106 31840 16140
rect 31930 16106 32098 16140
rect 32904 17584 32972 17618
rect 32904 17056 32972 17090
rect 33546 17588 33614 17622
rect 33546 16078 33614 16112
<< locali >>
rect 2376 26468 2472 26502
rect 3182 26468 3278 26502
rect 2376 26406 2410 26468
rect 1136 24868 1232 24902
rect 1942 24868 2038 24902
rect 1136 24806 1170 24868
rect 2004 24806 2038 24868
rect 1296 24766 1312 24800
rect 1350 24766 1366 24800
rect 1424 24766 1440 24800
rect 1478 24766 1494 24800
rect 1552 24766 1568 24800
rect 1606 24766 1622 24800
rect 1680 24766 1696 24800
rect 1734 24766 1750 24800
rect 1808 24766 1824 24800
rect 1862 24766 1878 24800
rect 1250 24707 1284 24723
rect 1250 23115 1284 23131
rect 1378 24707 1412 24723
rect 1378 23115 1412 23131
rect 1506 24707 1540 24723
rect 1506 23115 1540 23131
rect 1634 24707 1668 24723
rect 1634 23115 1668 23131
rect 1762 24707 1796 24723
rect 1762 23115 1796 23131
rect 1890 24707 1924 24723
rect 1890 23115 1924 23131
rect 1296 23038 1312 23072
rect 1350 23038 1366 23072
rect 1424 23038 1440 23072
rect 1478 23038 1494 23072
rect 1552 23038 1568 23072
rect 1606 23038 1622 23072
rect 1680 23038 1696 23072
rect 1734 23038 1750 23072
rect 1808 23038 1824 23072
rect 1862 23038 1878 23072
rect 1136 22970 1170 23032
rect 3244 26406 3278 26468
rect 2536 26366 2552 26400
rect 2590 26366 2606 26400
rect 2664 26366 2680 26400
rect 2718 26366 2734 26400
rect 2792 26366 2808 26400
rect 2846 26366 2862 26400
rect 2920 26366 2936 26400
rect 2974 26366 2990 26400
rect 3048 26366 3064 26400
rect 3102 26366 3118 26400
rect 2490 26307 2524 26323
rect 2490 24715 2524 24731
rect 2618 26307 2652 26323
rect 2618 24715 2652 24731
rect 2746 26307 2780 26323
rect 2746 24715 2780 24731
rect 2874 26307 2908 26323
rect 2874 24715 2908 24731
rect 3002 26307 3036 26323
rect 3002 24715 3036 24731
rect 3130 26307 3164 26323
rect 3130 24715 3164 24731
rect 2536 24638 2552 24672
rect 2590 24638 2606 24672
rect 2664 24638 2680 24672
rect 2718 24638 2734 24672
rect 2792 24638 2808 24672
rect 2846 24638 2862 24672
rect 2920 24638 2936 24672
rect 2974 24638 2990 24672
rect 3048 24638 3064 24672
rect 3102 24638 3118 24672
rect 2376 24570 2410 24632
rect 11516 26468 11612 26502
rect 12322 26468 12418 26502
rect 11516 26406 11550 26468
rect 3244 24570 3278 24632
rect 2376 24536 2472 24570
rect 3182 24536 3278 24570
rect 10276 24868 10372 24902
rect 11082 24868 11178 24902
rect 10276 24806 10310 24868
rect 2004 22970 2038 23032
rect 1136 22936 1232 22970
rect 1942 22936 2038 22970
rect 11144 24806 11178 24868
rect 10436 24766 10452 24800
rect 10490 24766 10506 24800
rect 10564 24766 10580 24800
rect 10618 24766 10634 24800
rect 10692 24766 10708 24800
rect 10746 24766 10762 24800
rect 10820 24766 10836 24800
rect 10874 24766 10890 24800
rect 10948 24766 10964 24800
rect 11002 24766 11018 24800
rect 10390 24707 10424 24723
rect 10390 23115 10424 23131
rect 10518 24707 10552 24723
rect 10518 23115 10552 23131
rect 10646 24707 10680 24723
rect 10646 23115 10680 23131
rect 10774 24707 10808 24723
rect 10774 23115 10808 23131
rect 10902 24707 10936 24723
rect 10902 23115 10936 23131
rect 11030 24707 11064 24723
rect 11030 23115 11064 23131
rect 10436 23038 10452 23072
rect 10490 23038 10506 23072
rect 10564 23038 10580 23072
rect 10618 23038 10634 23072
rect 10692 23038 10708 23072
rect 10746 23038 10762 23072
rect 10820 23038 10836 23072
rect 10874 23038 10890 23072
rect 10948 23038 10964 23072
rect 11002 23038 11018 23072
rect 10276 22970 10310 23032
rect 12384 26406 12418 26468
rect 11676 26366 11692 26400
rect 11730 26366 11746 26400
rect 11804 26366 11820 26400
rect 11858 26366 11874 26400
rect 11932 26366 11948 26400
rect 11986 26366 12002 26400
rect 12060 26366 12076 26400
rect 12114 26366 12130 26400
rect 12188 26366 12204 26400
rect 12242 26366 12258 26400
rect 11630 26307 11664 26323
rect 11630 24715 11664 24731
rect 11758 26307 11792 26323
rect 11758 24715 11792 24731
rect 11886 26307 11920 26323
rect 11886 24715 11920 24731
rect 12014 26307 12048 26323
rect 12014 24715 12048 24731
rect 12142 26307 12176 26323
rect 12142 24715 12176 24731
rect 12270 26307 12304 26323
rect 12270 24715 12304 24731
rect 11676 24638 11692 24672
rect 11730 24638 11746 24672
rect 11804 24638 11820 24672
rect 11858 24638 11874 24672
rect 11932 24638 11948 24672
rect 11986 24638 12002 24672
rect 12060 24638 12076 24672
rect 12114 24638 12130 24672
rect 12188 24638 12204 24672
rect 12242 24638 12258 24672
rect 11516 24570 11550 24632
rect 20706 26468 20802 26502
rect 21512 26468 21608 26502
rect 20706 26406 20740 26468
rect 12384 24570 12418 24632
rect 11516 24536 11612 24570
rect 12322 24536 12418 24570
rect 19466 24868 19562 24902
rect 20272 24868 20368 24902
rect 19466 24806 19500 24868
rect 11144 22970 11178 23032
rect 10276 22936 10372 22970
rect 11082 22936 11178 22970
rect 20334 24806 20368 24868
rect 19626 24766 19642 24800
rect 19680 24766 19696 24800
rect 19754 24766 19770 24800
rect 19808 24766 19824 24800
rect 19882 24766 19898 24800
rect 19936 24766 19952 24800
rect 20010 24766 20026 24800
rect 20064 24766 20080 24800
rect 20138 24766 20154 24800
rect 20192 24766 20208 24800
rect 19580 24707 19614 24723
rect 19580 23115 19614 23131
rect 19708 24707 19742 24723
rect 19708 23115 19742 23131
rect 19836 24707 19870 24723
rect 19836 23115 19870 23131
rect 19964 24707 19998 24723
rect 19964 23115 19998 23131
rect 20092 24707 20126 24723
rect 20092 23115 20126 23131
rect 20220 24707 20254 24723
rect 20220 23115 20254 23131
rect 19626 23038 19642 23072
rect 19680 23038 19696 23072
rect 19754 23038 19770 23072
rect 19808 23038 19824 23072
rect 19882 23038 19898 23072
rect 19936 23038 19952 23072
rect 20010 23038 20026 23072
rect 20064 23038 20080 23072
rect 20138 23038 20154 23072
rect 20192 23038 20208 23072
rect 19466 22970 19500 23032
rect 21574 26406 21608 26468
rect 20866 26366 20882 26400
rect 20920 26366 20936 26400
rect 20994 26366 21010 26400
rect 21048 26366 21064 26400
rect 21122 26366 21138 26400
rect 21176 26366 21192 26400
rect 21250 26366 21266 26400
rect 21304 26366 21320 26400
rect 21378 26366 21394 26400
rect 21432 26366 21448 26400
rect 20820 26307 20854 26323
rect 20820 24715 20854 24731
rect 20948 26307 20982 26323
rect 20948 24715 20982 24731
rect 21076 26307 21110 26323
rect 21076 24715 21110 24731
rect 21204 26307 21238 26323
rect 21204 24715 21238 24731
rect 21332 26307 21366 26323
rect 21332 24715 21366 24731
rect 21460 26307 21494 26323
rect 21460 24715 21494 24731
rect 20866 24638 20882 24672
rect 20920 24638 20936 24672
rect 20994 24638 21010 24672
rect 21048 24638 21064 24672
rect 21122 24638 21138 24672
rect 21176 24638 21192 24672
rect 21250 24638 21266 24672
rect 21304 24638 21320 24672
rect 21378 24638 21394 24672
rect 21432 24638 21448 24672
rect 20706 24570 20740 24632
rect 31215 25875 31311 25909
rect 33539 25875 33635 25909
rect 31215 25813 31249 25875
rect 33601 25813 33635 25875
rect 31421 25741 31437 25775
rect 33413 25741 33429 25775
rect 31353 25713 31387 25729
rect 31353 25629 31387 25645
rect 33463 25713 33497 25729
rect 33463 25629 33497 25645
rect 31421 25583 31437 25617
rect 33413 25583 33429 25617
rect 31215 25483 31249 25545
rect 33601 25483 33635 25545
rect 31215 25449 31311 25483
rect 33539 25449 33635 25483
rect 21574 24570 21608 24632
rect 20706 24536 20802 24570
rect 21512 24536 21608 24570
rect 20334 22970 20368 23032
rect 19466 22936 19562 22970
rect 20272 22936 20368 22970
rect 30220 20426 30316 20460
rect 32232 20426 32328 20460
rect 30220 20364 30254 20426
rect 32294 20364 32328 20426
rect 30400 20288 30416 20322
rect 30584 20288 30600 20322
rect 30658 20288 30674 20322
rect 30842 20288 30858 20322
rect 30916 20288 30932 20322
rect 31100 20288 31116 20322
rect 31174 20288 31190 20322
rect 31358 20288 31374 20322
rect 31432 20288 31448 20322
rect 31616 20288 31632 20322
rect 31690 20288 31706 20322
rect 31874 20288 31890 20322
rect 31948 20288 31964 20322
rect 32132 20288 32148 20322
rect 30354 20238 30388 20254
rect 30354 19646 30388 19662
rect 30612 20238 30646 20254
rect 30612 19646 30646 19662
rect 30870 20238 30904 20254
rect 30870 19646 30904 19662
rect 31128 20238 31162 20254
rect 31128 19646 31162 19662
rect 31386 20238 31420 20254
rect 31386 19646 31420 19662
rect 31644 20238 31678 20254
rect 31644 19646 31678 19662
rect 31902 20238 31936 20254
rect 31902 19646 31936 19662
rect 32160 20238 32194 20254
rect 32160 19646 32194 19662
rect 30400 19578 30416 19612
rect 30584 19578 30600 19612
rect 30658 19578 30674 19612
rect 30842 19578 30858 19612
rect 30916 19578 30932 19612
rect 31100 19578 31116 19612
rect 31174 19578 31190 19612
rect 31358 19578 31374 19612
rect 31432 19578 31448 19612
rect 31616 19578 31632 19612
rect 31690 19578 31706 19612
rect 31874 19578 31890 19612
rect 31948 19578 31964 19612
rect 32132 19578 32148 19612
rect 32294 19474 32328 19536
rect 30220 19440 30316 19474
rect 32232 19440 32328 19474
rect 33350 19626 33446 19660
rect 33714 19626 33810 19660
rect 33350 19564 33384 19626
rect 28638 19222 28734 19256
rect 32198 19222 32294 19256
rect 28638 19160 28672 19222
rect 32260 19160 32294 19222
rect 28818 19084 28834 19118
rect 29002 19084 29018 19118
rect 29076 19084 29092 19118
rect 29260 19084 29276 19118
rect 29334 19084 29350 19118
rect 29518 19084 29534 19118
rect 29592 19084 29608 19118
rect 29776 19084 29792 19118
rect 29850 19084 29866 19118
rect 30034 19084 30050 19118
rect 30108 19084 30124 19118
rect 30292 19084 30308 19118
rect 30366 19084 30382 19118
rect 30550 19084 30566 19118
rect 30624 19084 30640 19118
rect 30808 19084 30824 19118
rect 30882 19084 30898 19118
rect 31066 19084 31082 19118
rect 31140 19084 31156 19118
rect 31324 19084 31340 19118
rect 31398 19084 31414 19118
rect 31582 19084 31598 19118
rect 31656 19084 31672 19118
rect 31840 19084 31856 19118
rect 31914 19084 31930 19118
rect 32098 19084 32114 19118
rect 28772 19025 28806 19041
rect 28772 18433 28806 18449
rect 29030 19025 29064 19041
rect 29030 18433 29064 18449
rect 29288 19025 29322 19041
rect 29288 18433 29322 18449
rect 29546 19025 29580 19041
rect 29546 18433 29580 18449
rect 29804 19025 29838 19041
rect 29804 18433 29838 18449
rect 30062 19025 30096 19041
rect 30062 18433 30096 18449
rect 30320 19025 30354 19041
rect 30320 18433 30354 18449
rect 30578 19025 30612 19041
rect 30578 18433 30612 18449
rect 30836 19025 30870 19041
rect 30836 18433 30870 18449
rect 31094 19025 31128 19041
rect 31094 18433 31128 18449
rect 31352 19025 31386 19041
rect 31352 18433 31386 18449
rect 31610 19025 31644 19041
rect 31610 18433 31644 18449
rect 31868 19025 31902 19041
rect 31868 18433 31902 18449
rect 32126 19025 32160 19041
rect 32126 18433 32160 18449
rect 28818 18356 28834 18390
rect 29002 18356 29018 18390
rect 29076 18356 29092 18390
rect 29260 18356 29276 18390
rect 29334 18356 29350 18390
rect 29518 18356 29534 18390
rect 29592 18356 29608 18390
rect 29776 18356 29792 18390
rect 29850 18356 29866 18390
rect 30034 18356 30050 18390
rect 30108 18356 30124 18390
rect 30292 18356 30308 18390
rect 30366 18356 30382 18390
rect 30550 18356 30566 18390
rect 30624 18356 30640 18390
rect 30808 18356 30824 18390
rect 30882 18356 30898 18390
rect 31066 18356 31082 18390
rect 31140 18356 31156 18390
rect 31324 18356 31340 18390
rect 31398 18356 31414 18390
rect 31582 18356 31598 18390
rect 31656 18356 31672 18390
rect 31840 18356 31856 18390
rect 31914 18356 31930 18390
rect 32098 18356 32114 18390
rect 32260 18252 32294 18314
rect 28638 18218 28734 18252
rect 32198 18218 32294 18252
rect 32708 18642 32804 18676
rect 33072 18642 33168 18676
rect 32708 18580 32742 18642
rect 33134 18580 33168 18642
rect 32888 18504 32904 18538
rect 32972 18504 32988 18538
rect 29928 18102 30024 18136
rect 32198 18102 32294 18136
rect 29928 18040 29962 18102
rect 32260 18040 32294 18102
rect 30108 17964 30124 17998
rect 30292 17964 30308 17998
rect 30366 17964 30382 17998
rect 30550 17964 30566 17998
rect 30624 17964 30640 17998
rect 30808 17964 30824 17998
rect 30882 17964 30898 17998
rect 31066 17964 31082 17998
rect 31140 17964 31156 17998
rect 31324 17964 31340 17998
rect 31398 17964 31414 17998
rect 31582 17964 31598 17998
rect 31656 17964 31672 17998
rect 31840 17964 31856 17998
rect 31914 17964 31930 17998
rect 32098 17964 32114 17998
rect 30062 17905 30096 17921
rect 30062 17313 30096 17329
rect 30320 17905 30354 17921
rect 30320 17313 30354 17329
rect 30578 17905 30612 17921
rect 30578 17313 30612 17329
rect 30836 17905 30870 17921
rect 30836 17313 30870 17329
rect 31094 17905 31128 17921
rect 31094 17313 31128 17329
rect 31352 17905 31386 17921
rect 31352 17313 31386 17329
rect 31610 17905 31644 17921
rect 31610 17313 31644 17329
rect 31868 17905 31902 17921
rect 31868 17313 31902 17329
rect 32126 17905 32160 17921
rect 32126 17313 32160 17329
rect 30108 17236 30124 17270
rect 30292 17236 30308 17270
rect 30366 17236 30382 17270
rect 30550 17236 30566 17270
rect 30624 17236 30640 17270
rect 30808 17236 30824 17270
rect 30882 17236 30898 17270
rect 31066 17236 31082 17270
rect 31140 17236 31156 17270
rect 31324 17236 31340 17270
rect 31398 17236 31414 17270
rect 31582 17236 31598 17270
rect 31656 17236 31672 17270
rect 31840 17236 31856 17270
rect 31914 17236 31930 17270
rect 32098 17236 32114 17270
rect 32842 18445 32876 18461
rect 32842 18053 32876 18069
rect 33000 18445 33034 18461
rect 33000 18053 33034 18069
rect 32888 17976 32904 18010
rect 32972 17976 32988 18010
rect 32708 17872 32742 17934
rect 33134 17872 33168 17934
rect 32708 17838 32804 17872
rect 33072 17838 33168 17872
rect 33776 19564 33810 19626
rect 33530 19488 33546 19522
rect 33614 19488 33630 19522
rect 33484 19438 33518 19454
rect 33484 18046 33518 18062
rect 33642 19438 33676 19454
rect 33642 18046 33676 18062
rect 33530 17978 33546 18012
rect 33614 17978 33630 18012
rect 33350 17874 33384 17936
rect 33350 17840 33446 17874
rect 33714 17840 33810 17874
rect 32260 17132 32294 17194
rect 29928 17098 30024 17132
rect 32198 17098 32294 17132
rect 32708 17722 32804 17756
rect 33072 17722 33168 17756
rect 32708 17660 32742 17722
rect 33134 17660 33168 17722
rect 32888 17584 32904 17618
rect 32972 17584 32988 17618
rect 32842 17525 32876 17541
rect 32842 17133 32876 17149
rect 33000 17525 33034 17541
rect 33000 17133 33034 17149
rect 32888 17056 32904 17090
rect 32972 17056 32988 17090
rect 29928 16972 30024 17006
rect 32198 16972 32294 17006
rect 32260 16910 32294 16972
rect 32708 16952 32742 17014
rect 33134 16952 33168 17014
rect 32708 16918 32804 16952
rect 33072 16918 33168 16952
rect 33350 17726 33446 17760
rect 33714 17726 33810 17760
rect 33350 17664 33384 17726
rect 30108 16834 30124 16868
rect 30292 16834 30308 16868
rect 30366 16834 30382 16868
rect 30550 16834 30566 16868
rect 30624 16834 30640 16868
rect 30808 16834 30824 16868
rect 30882 16834 30898 16868
rect 31066 16834 31082 16868
rect 31140 16834 31156 16868
rect 31324 16834 31340 16868
rect 31398 16834 31414 16868
rect 31582 16834 31598 16868
rect 31656 16834 31672 16868
rect 31840 16834 31856 16868
rect 31914 16834 31930 16868
rect 32098 16834 32114 16868
rect 30062 16775 30096 16791
rect 30062 16183 30096 16199
rect 30320 16775 30354 16791
rect 30320 16183 30354 16199
rect 30578 16775 30612 16791
rect 30578 16183 30612 16199
rect 30836 16775 30870 16791
rect 30836 16183 30870 16199
rect 31094 16775 31128 16791
rect 31094 16183 31128 16199
rect 31352 16775 31386 16791
rect 31352 16183 31386 16199
rect 31610 16775 31644 16791
rect 31610 16183 31644 16199
rect 31868 16775 31902 16791
rect 31868 16183 31902 16199
rect 32126 16775 32160 16791
rect 32126 16183 32160 16199
rect 30108 16106 30124 16140
rect 30292 16106 30308 16140
rect 30366 16106 30382 16140
rect 30550 16106 30566 16140
rect 30624 16106 30640 16140
rect 30808 16106 30824 16140
rect 30882 16106 30898 16140
rect 31066 16106 31082 16140
rect 31140 16106 31156 16140
rect 31324 16106 31340 16140
rect 31398 16106 31414 16140
rect 31582 16106 31598 16140
rect 31656 16106 31672 16140
rect 31840 16106 31856 16140
rect 31914 16106 31930 16140
rect 32098 16106 32114 16140
rect 29928 16002 29962 16064
rect 32260 16002 32294 16064
rect 29928 15968 30024 16002
rect 32198 15968 32294 16002
rect 33530 17588 33546 17622
rect 33614 17588 33630 17622
rect 33484 17538 33518 17554
rect 33484 16146 33518 16162
rect 33642 17538 33676 17554
rect 33642 16146 33676 16162
rect 33530 16078 33546 16112
rect 33614 16078 33630 16112
rect 33350 15974 33384 16036
rect 33776 15974 33810 16036
rect 33350 15940 33446 15974
rect 33714 15940 33810 15974
<< viali >>
rect 2619 26468 3035 26502
rect 1379 24868 1795 24902
rect 1312 24766 1350 24800
rect 1440 24766 1478 24800
rect 1568 24766 1606 24800
rect 1696 24766 1734 24800
rect 1824 24766 1862 24800
rect 1250 24060 1284 24690
rect 1378 23148 1412 23778
rect 1506 24060 1540 24690
rect 1634 23148 1668 23778
rect 1762 24060 1796 24690
rect 1890 23148 1924 23778
rect 1312 23038 1350 23072
rect 1440 23038 1478 23072
rect 1568 23038 1606 23072
rect 1696 23038 1734 23072
rect 1824 23038 1862 23072
rect 2552 26366 2590 26400
rect 2680 26366 2718 26400
rect 2808 26366 2846 26400
rect 2936 26366 2974 26400
rect 3064 26366 3102 26400
rect 2490 25660 2524 26290
rect 2618 24748 2652 25378
rect 2746 25660 2780 26290
rect 2874 24748 2908 25378
rect 3002 25660 3036 26290
rect 3130 24748 3164 25378
rect 2552 24638 2590 24672
rect 2680 24638 2718 24672
rect 2808 24638 2846 24672
rect 2936 24638 2974 24672
rect 3064 24638 3102 24672
rect 11759 26468 12175 26502
rect 10519 24868 10935 24902
rect 10452 24766 10490 24800
rect 10580 24766 10618 24800
rect 10708 24766 10746 24800
rect 10836 24766 10874 24800
rect 10964 24766 11002 24800
rect 10390 24060 10424 24690
rect 10518 23148 10552 23778
rect 10646 24060 10680 24690
rect 10774 23148 10808 23778
rect 10902 24060 10936 24690
rect 11030 23148 11064 23778
rect 10452 23038 10490 23072
rect 10580 23038 10618 23072
rect 10708 23038 10746 23072
rect 10836 23038 10874 23072
rect 10964 23038 11002 23072
rect 11692 26366 11730 26400
rect 11820 26366 11858 26400
rect 11948 26366 11986 26400
rect 12076 26366 12114 26400
rect 12204 26366 12242 26400
rect 11630 25660 11664 26290
rect 11758 24748 11792 25378
rect 11886 25660 11920 26290
rect 12014 24748 12048 25378
rect 12142 25660 12176 26290
rect 12270 24748 12304 25378
rect 11692 24638 11730 24672
rect 11820 24638 11858 24672
rect 11948 24638 11986 24672
rect 12076 24638 12114 24672
rect 12204 24638 12242 24672
rect 20949 26468 21365 26502
rect 19709 24868 20125 24902
rect 19642 24766 19680 24800
rect 19770 24766 19808 24800
rect 19898 24766 19936 24800
rect 20026 24766 20064 24800
rect 20154 24766 20192 24800
rect 19580 24060 19614 24690
rect 19708 23148 19742 23778
rect 19836 24060 19870 24690
rect 19964 23148 19998 23778
rect 20092 24060 20126 24690
rect 20220 23148 20254 23778
rect 19642 23038 19680 23072
rect 19770 23038 19808 23072
rect 19898 23038 19936 23072
rect 20026 23038 20064 23072
rect 20154 23038 20192 23072
rect 20882 26366 20920 26400
rect 21010 26366 21048 26400
rect 21138 26366 21176 26400
rect 21266 26366 21304 26400
rect 21394 26366 21432 26400
rect 20820 25660 20854 26290
rect 20948 24748 20982 25378
rect 21076 25660 21110 26290
rect 21204 24748 21238 25378
rect 21332 25660 21366 26290
rect 21460 24748 21494 25378
rect 20882 24638 20920 24672
rect 21010 24638 21048 24672
rect 21138 24638 21176 24672
rect 21266 24638 21304 24672
rect 21394 24638 21432 24672
rect 33001 25741 33396 25775
rect 31353 25645 31387 25713
rect 33463 25645 33497 25713
rect 31454 25583 31849 25617
rect 32249 25449 32601 25483
rect 30416 20288 30584 20322
rect 30674 20288 30842 20322
rect 30932 20288 31100 20322
rect 31190 20288 31358 20322
rect 31448 20288 31616 20322
rect 31706 20288 31874 20322
rect 31964 20288 32132 20322
rect 30220 19536 30254 19950
rect 30354 19991 30388 20221
rect 30612 19679 30646 19909
rect 30870 19991 30904 20221
rect 31128 19679 31162 19909
rect 31386 19991 31420 20221
rect 31644 19679 31678 19909
rect 31902 19991 31936 20221
rect 32160 19679 32194 19909
rect 30416 19578 30584 19612
rect 30674 19578 30842 19612
rect 30932 19578 31100 19612
rect 31190 19578 31358 19612
rect 31448 19578 31616 19612
rect 31706 19578 31874 19612
rect 31964 19578 32132 19612
rect 30220 19474 30254 19536
rect 28834 19084 29002 19118
rect 29092 19084 29260 19118
rect 29350 19084 29518 19118
rect 29608 19084 29776 19118
rect 29866 19084 30034 19118
rect 30124 19084 30292 19118
rect 30382 19084 30550 19118
rect 30640 19084 30808 19118
rect 30898 19084 31066 19118
rect 31156 19084 31324 19118
rect 31414 19084 31582 19118
rect 31672 19084 31840 19118
rect 31930 19084 32098 19118
rect 28638 18314 28672 18737
rect 28772 18778 28806 19008
rect 29030 18466 29064 18696
rect 29288 18778 29322 19008
rect 29546 18466 29580 18696
rect 29804 18778 29838 19008
rect 30062 18466 30096 18696
rect 30320 18778 30354 19008
rect 30578 18466 30612 18696
rect 30836 18778 30870 19008
rect 31094 18466 31128 18696
rect 31352 18778 31386 19008
rect 31610 18466 31644 18696
rect 31868 18778 31902 19008
rect 32126 18466 32160 18696
rect 28834 18356 29002 18390
rect 29092 18356 29260 18390
rect 29350 18356 29518 18390
rect 29608 18356 29776 18390
rect 29866 18356 30034 18390
rect 30124 18356 30292 18390
rect 30382 18356 30550 18390
rect 30640 18356 30808 18390
rect 30898 18356 31066 18390
rect 31156 18356 31324 18390
rect 31414 18356 31582 18390
rect 31672 18356 31840 18390
rect 31930 18356 32098 18390
rect 28638 18252 28672 18314
rect 32904 18504 32972 18538
rect 32708 18199 32742 18315
rect 30124 17964 30292 17998
rect 30382 17964 30550 17998
rect 30640 17964 30808 17998
rect 30898 17964 31066 17998
rect 31156 17964 31324 17998
rect 31414 17964 31582 17998
rect 31672 17964 31840 17998
rect 31930 17964 32098 17998
rect 29928 17194 29962 17617
rect 30062 17658 30096 17888
rect 30320 17346 30354 17576
rect 30578 17658 30612 17888
rect 30836 17346 30870 17576
rect 31094 17658 31128 17888
rect 31352 17346 31386 17576
rect 31610 17658 31644 17888
rect 31868 17346 31902 17576
rect 32126 17658 32160 17888
rect 30124 17236 30292 17270
rect 30382 17236 30550 17270
rect 30640 17236 30808 17270
rect 30898 17236 31066 17270
rect 31156 17236 31324 17270
rect 31414 17236 31582 17270
rect 31672 17236 31840 17270
rect 31930 17236 32098 17270
rect 29928 17132 29962 17194
rect 32842 18069 32876 18445
rect 33000 18069 33034 18445
rect 32904 17976 32972 18010
rect 33546 19488 33614 19522
rect 33484 18079 33518 18492
rect 33642 18079 33676 18492
rect 33546 17978 33614 18012
rect 33776 17936 33810 18400
rect 33776 17874 33810 17936
rect 32904 17584 32972 17618
rect 32708 17279 32742 17395
rect 32842 17149 32876 17525
rect 33000 17149 33034 17525
rect 32904 17056 32972 17090
rect 29928 16910 29962 16972
rect 29928 16487 29962 16910
rect 30124 16834 30292 16868
rect 30382 16834 30550 16868
rect 30640 16834 30808 16868
rect 30898 16834 31066 16868
rect 31156 16834 31324 16868
rect 31414 16834 31582 16868
rect 31672 16834 31840 16868
rect 31930 16834 32098 16868
rect 30062 16528 30096 16758
rect 30320 16216 30354 16446
rect 30578 16528 30612 16758
rect 30836 16216 30870 16446
rect 31094 16528 31128 16758
rect 31352 16216 31386 16446
rect 31610 16528 31644 16758
rect 31868 16216 31902 16446
rect 32126 16528 32160 16758
rect 30124 16106 30292 16140
rect 30382 16106 30550 16140
rect 30640 16106 30808 16140
rect 30898 16106 31066 16140
rect 31156 16106 31324 16140
rect 31414 16106 31582 16140
rect 31672 16106 31840 16140
rect 31930 16106 32098 16140
rect 33776 17664 33810 17726
rect 33546 17588 33614 17622
rect 33484 17108 33518 17521
rect 33642 17108 33676 17521
rect 33776 17200 33810 17664
rect 33546 16078 33614 16112
<< metal1 >>
rect 770 33300 1200 33320
rect 10140 33300 10340 33320
rect 19330 33300 19530 33320
rect 770 33140 19530 33300
rect 770 33120 1200 33140
rect 1000 33100 1200 33120
rect 1000 32980 1040 33100
rect 1160 32980 1200 33100
rect 1000 32940 1200 32980
rect 10140 33100 10340 33140
rect 10140 32980 10180 33100
rect 10300 32980 10340 33100
rect 10140 32940 10340 32980
rect 19330 33100 19530 33140
rect 19330 32980 19370 33100
rect 19490 32980 19530 33100
rect 19330 32940 19530 32980
rect 2600 26502 3060 26540
rect 2600 26468 2619 26502
rect 3035 26468 3060 26502
rect 2600 26420 3060 26468
rect 11740 26502 12200 26540
rect 11740 26468 11759 26502
rect 12175 26468 12200 26502
rect 11740 26420 12200 26468
rect 20930 26502 21390 26540
rect 20930 26468 20949 26502
rect 21365 26468 21390 26502
rect 20930 26420 21390 26468
rect 2480 26400 3180 26420
rect 2480 26366 2552 26400
rect 2590 26366 2680 26400
rect 2718 26366 2808 26400
rect 2846 26366 2936 26400
rect 2974 26366 3064 26400
rect 3102 26366 3180 26400
rect 2480 26290 3180 26366
rect 1580 26060 1740 26080
rect 1580 25940 1600 26060
rect 1720 25940 1740 26060
rect 1580 25140 1740 25940
rect 2480 25660 2490 26290
rect 2524 25660 2746 26290
rect 2780 25660 3002 26290
rect 3036 26240 3180 26290
rect 11620 26400 12320 26420
rect 11620 26366 11692 26400
rect 11730 26366 11820 26400
rect 11858 26366 11948 26400
rect 11986 26366 12076 26400
rect 12114 26366 12204 26400
rect 12242 26366 12320 26400
rect 11620 26290 12320 26366
rect 3036 26220 4300 26240
rect 3036 26060 4120 26220
rect 4280 26060 4300 26220
rect 9900 26200 10100 26240
rect 9640 26180 10100 26200
rect 9640 26080 9660 26180
rect 9780 26080 10100 26180
rect 9640 26060 10100 26080
rect 3036 26040 4300 26060
rect 9900 26040 10100 26060
rect 10720 26060 10880 26080
rect 3036 25660 3180 26040
rect 2480 25640 3180 25660
rect 2612 25378 2658 25390
rect 2612 25140 2618 25378
rect 1500 24940 2618 25140
rect 1360 24902 1820 24940
rect 1360 24868 1379 24902
rect 1795 24868 1820 24902
rect 1360 24820 1820 24868
rect 1240 24800 1940 24820
rect 1240 24766 1312 24800
rect 1350 24766 1440 24800
rect 1478 24766 1568 24800
rect 1606 24766 1696 24800
rect 1734 24766 1824 24800
rect 1862 24766 1940 24800
rect 1240 24690 1940 24766
rect 2612 24748 2618 24940
rect 2652 25140 2658 25378
rect 2868 25378 2914 25390
rect 2868 25140 2874 25378
rect 2652 24940 2874 25140
rect 2652 24748 2658 24940
rect 2612 24736 2658 24748
rect 2868 24748 2874 24940
rect 2908 25140 2914 25378
rect 3124 25378 3170 25390
rect 3124 25140 3130 25378
rect 2908 24940 3130 25140
rect 2908 24748 2914 24940
rect 2868 24736 2914 24748
rect 3124 24748 3130 24940
rect 3164 25140 3170 25378
rect 3164 24940 3180 25140
rect 3164 24748 3170 24940
rect 3124 24736 3170 24748
rect 1240 24060 1250 24690
rect 1284 24060 1506 24690
rect 1540 24060 1762 24690
rect 1796 24060 1940 24690
rect 2540 24672 3120 24680
rect 2540 24638 2552 24672
rect 2590 24638 2680 24672
rect 2718 24638 2808 24672
rect 2846 24638 2936 24672
rect 2974 24638 3064 24672
rect 3102 24638 3120 24672
rect 2540 24620 3120 24638
rect 1244 24048 1290 24060
rect 1500 24048 1546 24060
rect 1756 24048 1802 24060
rect 1372 23778 1418 23790
rect 1372 23440 1378 23778
rect 1360 23240 1378 23440
rect 1372 23148 1378 23240
rect 1412 23440 1418 23778
rect 1628 23778 1674 23790
rect 1628 23440 1634 23778
rect 1412 23240 1634 23440
rect 1412 23148 1418 23240
rect 1372 23136 1418 23148
rect 1628 23148 1634 23240
rect 1668 23440 1674 23778
rect 1884 23778 1930 23790
rect 1884 23440 1890 23778
rect 1668 23240 1890 23440
rect 1668 23148 1674 23240
rect 1628 23136 1674 23148
rect 1884 23148 1890 23240
rect 1924 23440 1930 23778
rect 1924 23240 2180 23440
rect 1924 23148 1930 23240
rect 1884 23136 1930 23148
rect 1280 23072 1880 23080
rect 1280 23038 1312 23072
rect 1350 23038 1440 23072
rect 1478 23038 1568 23072
rect 1606 23038 1696 23072
rect 1734 23038 1824 23072
rect 1862 23038 1880 23072
rect 1280 23020 1880 23038
rect 1980 22880 2180 23240
rect 770 22860 3700 22880
rect 770 22700 3520 22860
rect 3680 22700 3700 22860
rect 9920 22860 10080 26040
rect 10720 25940 10740 26060
rect 10860 25940 10880 26060
rect 10720 25140 10880 25940
rect 11620 25660 11630 26290
rect 11664 25660 11886 26290
rect 11920 25660 12142 26290
rect 12176 26240 12320 26290
rect 20810 26400 21510 26420
rect 20810 26366 20882 26400
rect 20920 26366 21010 26400
rect 21048 26366 21138 26400
rect 21176 26366 21266 26400
rect 21304 26366 21394 26400
rect 21432 26366 21510 26400
rect 20810 26290 21510 26366
rect 12176 26220 13440 26240
rect 12176 26060 13260 26220
rect 13420 26060 13440 26220
rect 19040 26200 19240 26240
rect 18780 26180 19240 26200
rect 18780 26080 18800 26180
rect 18920 26080 19240 26180
rect 18780 26060 19240 26080
rect 12176 26040 13440 26060
rect 19040 26040 19240 26060
rect 19910 26060 20070 26080
rect 12176 25660 12320 26040
rect 11620 25640 12320 25660
rect 11752 25378 11798 25390
rect 11752 25140 11758 25378
rect 10640 24940 11758 25140
rect 10500 24902 10960 24940
rect 10500 24868 10519 24902
rect 10935 24868 10960 24902
rect 10500 24820 10960 24868
rect 10380 24800 11080 24820
rect 10380 24766 10452 24800
rect 10490 24766 10580 24800
rect 10618 24766 10708 24800
rect 10746 24766 10836 24800
rect 10874 24766 10964 24800
rect 11002 24766 11080 24800
rect 10380 24690 11080 24766
rect 11752 24748 11758 24940
rect 11792 25140 11798 25378
rect 12008 25378 12054 25390
rect 12008 25140 12014 25378
rect 11792 24940 12014 25140
rect 11792 24748 11798 24940
rect 11752 24736 11798 24748
rect 12008 24748 12014 24940
rect 12048 25140 12054 25378
rect 12264 25378 12310 25390
rect 12264 25140 12270 25378
rect 12048 24940 12270 25140
rect 12048 24748 12054 24940
rect 12008 24736 12054 24748
rect 12264 24748 12270 24940
rect 12304 25140 12310 25378
rect 12304 24940 12320 25140
rect 12304 24748 12310 24940
rect 12264 24736 12310 24748
rect 10380 24060 10390 24690
rect 10424 24060 10646 24690
rect 10680 24060 10902 24690
rect 10936 24060 11080 24690
rect 11680 24672 12260 24680
rect 11680 24638 11692 24672
rect 11730 24638 11820 24672
rect 11858 24638 11948 24672
rect 11986 24638 12076 24672
rect 12114 24638 12204 24672
rect 12242 24638 12260 24672
rect 11680 24620 12260 24638
rect 10384 24048 10430 24060
rect 10640 24048 10686 24060
rect 10896 24048 10942 24060
rect 10512 23778 10558 23790
rect 10512 23440 10518 23778
rect 10500 23240 10518 23440
rect 10512 23148 10518 23240
rect 10552 23440 10558 23778
rect 10768 23778 10814 23790
rect 10768 23440 10774 23778
rect 10552 23240 10774 23440
rect 10552 23148 10558 23240
rect 10512 23136 10558 23148
rect 10768 23148 10774 23240
rect 10808 23440 10814 23778
rect 11024 23778 11070 23790
rect 11024 23440 11030 23778
rect 10808 23240 11030 23440
rect 10808 23148 10814 23240
rect 10768 23136 10814 23148
rect 11024 23148 11030 23240
rect 11064 23440 11070 23778
rect 11064 23240 11320 23440
rect 11064 23148 11070 23240
rect 11024 23136 11070 23148
rect 10420 23072 11020 23080
rect 10420 23038 10452 23072
rect 10490 23038 10580 23072
rect 10618 23038 10708 23072
rect 10746 23038 10836 23072
rect 10874 23038 10964 23072
rect 11002 23038 11020 23072
rect 10420 23020 11020 23038
rect 11120 22880 11320 23240
rect 10140 22860 12840 22880
rect 9920 22700 12660 22860
rect 12820 22700 12840 22860
rect 19060 22860 19220 26040
rect 19910 25940 19930 26060
rect 20050 25940 20070 26060
rect 19910 25140 20070 25940
rect 20810 25660 20820 26290
rect 20854 25660 21076 26290
rect 21110 25660 21332 26290
rect 21366 26240 21510 26290
rect 21366 26220 22630 26240
rect 21366 26060 22450 26220
rect 22610 26060 22630 26220
rect 28230 26220 28660 26240
rect 34330 26220 34760 26240
rect 28230 26200 31700 26220
rect 27970 26180 31700 26200
rect 27970 26080 27990 26180
rect 28110 26080 31700 26180
rect 27970 26060 31700 26080
rect 21366 26040 22630 26060
rect 28230 26040 28660 26060
rect 21366 25660 21510 26040
rect 20810 25640 21510 25660
rect 20942 25378 20988 25390
rect 20942 25140 20948 25378
rect 19830 24940 20948 25140
rect 19690 24902 20150 24940
rect 19690 24868 19709 24902
rect 20125 24868 20150 24902
rect 19690 24820 20150 24868
rect 19570 24800 20270 24820
rect 19570 24766 19642 24800
rect 19680 24766 19770 24800
rect 19808 24766 19898 24800
rect 19936 24766 20026 24800
rect 20064 24766 20154 24800
rect 20192 24766 20270 24800
rect 19570 24690 20270 24766
rect 20942 24748 20948 24940
rect 20982 25140 20988 25378
rect 21198 25378 21244 25390
rect 21198 25140 21204 25378
rect 20982 24940 21204 25140
rect 20982 24748 20988 24940
rect 20942 24736 20988 24748
rect 21198 24748 21204 24940
rect 21238 25140 21244 25378
rect 21454 25378 21500 25390
rect 21454 25140 21460 25378
rect 21238 24940 21460 25140
rect 21238 24748 21244 24940
rect 21198 24736 21244 24748
rect 21454 24748 21460 24940
rect 21494 25140 21500 25378
rect 21494 24940 21510 25140
rect 21494 24748 21500 24940
rect 21454 24736 21500 24748
rect 19570 24060 19580 24690
rect 19614 24060 19836 24690
rect 19870 24060 20092 24690
rect 20126 24060 20270 24690
rect 20870 24672 21450 24680
rect 20870 24638 20882 24672
rect 20920 24638 21010 24672
rect 21048 24638 21138 24672
rect 21176 24638 21266 24672
rect 21304 24638 21394 24672
rect 21432 24638 21450 24672
rect 20870 24620 21450 24638
rect 19574 24048 19620 24060
rect 19830 24048 19876 24060
rect 20086 24048 20132 24060
rect 19702 23778 19748 23790
rect 19702 23440 19708 23778
rect 19690 23240 19708 23440
rect 19702 23148 19708 23240
rect 19742 23440 19748 23778
rect 19958 23778 20004 23790
rect 19958 23440 19964 23778
rect 19742 23240 19964 23440
rect 19742 23148 19748 23240
rect 19702 23136 19748 23148
rect 19958 23148 19964 23240
rect 19998 23440 20004 23778
rect 20214 23778 20260 23790
rect 20214 23440 20220 23778
rect 19998 23240 20220 23440
rect 19998 23148 20004 23240
rect 19958 23136 20004 23148
rect 20214 23148 20220 23240
rect 20254 23440 20260 23778
rect 20254 23240 20510 23440
rect 20254 23148 20260 23240
rect 20214 23136 20260 23148
rect 19610 23072 20210 23080
rect 19610 23038 19642 23072
rect 19680 23038 19770 23072
rect 19808 23038 19898 23072
rect 19936 23038 20026 23072
rect 20064 23038 20154 23072
rect 20192 23038 20210 23072
rect 19610 23020 20210 23038
rect 20310 22880 20510 23240
rect 28480 23150 28640 26040
rect 31347 25713 31393 25725
rect 31347 25645 31353 25713
rect 31387 25645 31393 25713
rect 31347 25633 31393 25645
rect 31550 25623 31700 26060
rect 33120 26200 34760 26220
rect 33120 26080 33890 26200
rect 34010 26080 34760 26200
rect 33120 26060 34760 26080
rect 33120 25781 33270 26060
rect 34330 26040 34760 26060
rect 32989 25775 33408 25781
rect 32989 25741 33001 25775
rect 33396 25741 33408 25775
rect 32989 25735 33408 25741
rect 33120 25730 33270 25735
rect 33460 25725 34030 25730
rect 33457 25713 34030 25725
rect 33457 25645 33463 25713
rect 33497 25645 34030 25713
rect 33457 25633 34030 25645
rect 33460 25630 34030 25633
rect 31442 25617 31861 25623
rect 31442 25583 31454 25617
rect 31849 25583 31861 25617
rect 31442 25577 31861 25583
rect 32360 25489 32490 25490
rect 32237 25483 32613 25489
rect 32237 25449 32249 25483
rect 32601 25449 32613 25483
rect 32237 25443 32613 25449
rect 32360 25410 32490 25443
rect 32360 25320 32380 25410
rect 32470 25320 32490 25410
rect 32360 25300 32490 25320
rect 28480 23030 28500 23150
rect 28620 23030 28640 23150
rect 28480 23010 28640 23030
rect 19330 22860 22030 22880
rect 19060 22700 21850 22860
rect 22010 22700 22030 22860
rect 770 22680 3700 22700
rect 10140 22680 12840 22700
rect 19330 22680 22030 22700
rect 3310 22260 3500 22680
rect 3310 22240 12830 22260
rect 3310 22080 12660 22240
rect 12810 22080 12830 22240
rect 3310 22060 12830 22080
rect 21810 22240 28890 22260
rect 21810 22080 21830 22240
rect 22010 22080 28720 22240
rect 28870 22080 28890 22240
rect 21810 22060 28890 22080
rect 30404 20322 30596 20328
rect 30404 20288 30416 20322
rect 30584 20288 30596 20322
rect 30404 20282 30596 20288
rect 30662 20322 30854 20328
rect 30662 20288 30674 20322
rect 30842 20288 30854 20322
rect 30662 20282 30854 20288
rect 30920 20322 31112 20328
rect 30920 20288 30932 20322
rect 31100 20288 31112 20322
rect 30920 20282 31112 20288
rect 31178 20322 31370 20328
rect 31178 20288 31190 20322
rect 31358 20288 31370 20322
rect 31178 20282 31370 20288
rect 31436 20322 31628 20328
rect 31436 20288 31448 20322
rect 31616 20288 31628 20322
rect 31436 20282 31628 20288
rect 31694 20322 31886 20328
rect 31694 20288 31706 20322
rect 31874 20288 31886 20322
rect 31694 20282 31886 20288
rect 31952 20322 32144 20328
rect 31952 20288 31964 20322
rect 32132 20288 32144 20322
rect 31952 20282 32144 20288
rect 30348 20221 30394 20233
rect 30348 20180 30354 20221
rect 28480 20030 30354 20180
rect 28480 18970 28640 20030
rect 30348 19991 30354 20030
rect 30388 20180 30394 20221
rect 30864 20221 30910 20233
rect 30864 20180 30870 20221
rect 30388 20030 30870 20180
rect 30388 19991 30394 20030
rect 30348 19979 30394 19991
rect 30864 19991 30870 20030
rect 30904 20180 30910 20221
rect 31380 20221 31426 20233
rect 31380 20180 31386 20221
rect 30904 20030 31386 20180
rect 30904 19991 30910 20030
rect 30864 19979 30910 19991
rect 31380 19991 31386 20030
rect 31420 20180 31426 20221
rect 31896 20221 31942 20233
rect 31896 20180 31902 20221
rect 31420 20030 31902 20180
rect 31420 19991 31426 20030
rect 31380 19979 31426 19991
rect 31896 19991 31902 20030
rect 31936 20180 31942 20221
rect 33870 20210 34030 25630
rect 33850 20180 34050 20210
rect 31936 20160 34050 20180
rect 31936 20050 33690 20160
rect 33790 20050 34050 20160
rect 31936 20030 34050 20050
rect 31936 19991 31942 20030
rect 33850 20010 34050 20030
rect 31896 19979 31942 19991
rect 30214 19950 30260 19962
rect 30214 19870 30220 19950
rect 30210 19720 30220 19870
rect 30214 19474 30220 19720
rect 30254 19870 30260 19950
rect 30606 19909 30652 19921
rect 30606 19870 30612 19909
rect 30254 19720 30612 19870
rect 30254 19474 30260 19720
rect 30606 19679 30612 19720
rect 30646 19870 30652 19909
rect 31122 19909 31168 19921
rect 31122 19870 31128 19909
rect 30646 19720 31128 19870
rect 30646 19679 30652 19720
rect 30606 19667 30652 19679
rect 31122 19679 31128 19720
rect 31162 19870 31168 19909
rect 31638 19909 31684 19921
rect 31638 19870 31644 19909
rect 31162 19720 31644 19870
rect 31162 19679 31168 19720
rect 31122 19667 31168 19679
rect 31638 19679 31644 19720
rect 31678 19870 31684 19909
rect 32154 19909 32200 19921
rect 32154 19870 32160 19909
rect 31678 19720 32160 19870
rect 31678 19679 31684 19720
rect 31638 19667 31684 19679
rect 32154 19679 32160 19720
rect 32194 19870 32200 19909
rect 32194 19850 34030 19870
rect 32194 19740 33890 19850
rect 34010 19740 34030 19850
rect 32194 19720 34030 19740
rect 32194 19679 32200 19720
rect 32154 19667 32200 19679
rect 32790 19620 32800 19630
rect 30400 19612 32800 19620
rect 30400 19578 30416 19612
rect 30584 19578 30674 19612
rect 30842 19578 30932 19612
rect 31100 19578 31190 19612
rect 31358 19578 31448 19612
rect 31616 19578 31706 19612
rect 31874 19578 31964 19612
rect 32132 19578 32800 19612
rect 30400 19550 32800 19578
rect 32790 19540 32800 19550
rect 32890 19540 32900 19630
rect 33534 19522 33626 19528
rect 33534 19488 33546 19522
rect 33614 19488 33626 19522
rect 33534 19482 33626 19488
rect 30214 19462 30260 19474
rect 28822 19118 29014 19124
rect 28822 19084 28834 19118
rect 29002 19084 29014 19118
rect 28822 19078 29014 19084
rect 29080 19118 29272 19124
rect 29080 19084 29092 19118
rect 29260 19084 29272 19118
rect 29080 19078 29272 19084
rect 29338 19118 29530 19124
rect 29338 19084 29350 19118
rect 29518 19084 29530 19118
rect 29338 19078 29530 19084
rect 29596 19118 29788 19124
rect 29596 19084 29608 19118
rect 29776 19084 29788 19118
rect 29596 19078 29788 19084
rect 29854 19118 30046 19124
rect 29854 19084 29866 19118
rect 30034 19084 30046 19118
rect 29854 19078 30046 19084
rect 30112 19118 30304 19124
rect 30112 19084 30124 19118
rect 30292 19084 30304 19118
rect 30112 19078 30304 19084
rect 30370 19118 30562 19124
rect 30370 19084 30382 19118
rect 30550 19084 30562 19118
rect 30370 19078 30562 19084
rect 30628 19118 30820 19124
rect 30628 19084 30640 19118
rect 30808 19084 30820 19118
rect 30628 19078 30820 19084
rect 30886 19118 31078 19124
rect 30886 19084 30898 19118
rect 31066 19084 31078 19118
rect 30886 19078 31078 19084
rect 31144 19118 31336 19124
rect 31144 19084 31156 19118
rect 31324 19084 31336 19118
rect 31144 19078 31336 19084
rect 31402 19118 31594 19124
rect 31402 19084 31414 19118
rect 31582 19084 31594 19118
rect 31402 19078 31594 19084
rect 31660 19118 31852 19124
rect 31660 19084 31672 19118
rect 31840 19084 31852 19118
rect 31660 19078 31852 19084
rect 31918 19118 32110 19124
rect 31918 19084 31930 19118
rect 32098 19084 32110 19118
rect 31918 19078 32110 19084
rect 28766 19008 28812 19020
rect 28766 18970 28772 19008
rect 28480 18820 28772 18970
rect 28766 18778 28772 18820
rect 28806 18970 28812 19008
rect 29282 19008 29328 19020
rect 29282 18970 29288 19008
rect 28806 18820 29288 18970
rect 28806 18778 28812 18820
rect 28766 18766 28812 18778
rect 29282 18778 29288 18820
rect 29322 18970 29328 19008
rect 29798 19008 29844 19020
rect 29798 18970 29804 19008
rect 29322 18820 29804 18970
rect 29322 18778 29328 18820
rect 29282 18766 29328 18778
rect 29798 18778 29804 18820
rect 29838 18970 29844 19008
rect 30314 19008 30360 19020
rect 30314 18970 30320 19008
rect 29838 18820 30320 18970
rect 29838 18778 29844 18820
rect 29798 18766 29844 18778
rect 30314 18778 30320 18820
rect 30354 18970 30360 19008
rect 30830 19008 30876 19020
rect 30830 18970 30836 19008
rect 30354 18820 30836 18970
rect 30354 18778 30360 18820
rect 30314 18766 30360 18778
rect 30830 18778 30836 18820
rect 30870 18970 30876 19008
rect 31346 19008 31392 19020
rect 31346 18970 31352 19008
rect 30870 18820 31352 18970
rect 30870 18778 30876 18820
rect 30830 18766 30876 18778
rect 31346 18778 31352 18820
rect 31386 18970 31392 19008
rect 31862 19008 31908 19020
rect 31862 18970 31868 19008
rect 31386 18820 31868 18970
rect 31386 18778 31392 18820
rect 31346 18766 31392 18778
rect 31862 18778 31868 18820
rect 31902 18970 31908 19008
rect 31902 18820 31910 18970
rect 33850 18890 34050 18910
rect 34300 18890 34730 18910
rect 33850 18860 34730 18890
rect 31902 18778 31908 18820
rect 31862 18766 31908 18778
rect 32890 18760 34730 18860
rect 28632 18737 28678 18749
rect 28632 18650 28638 18737
rect 28480 18252 28638 18650
rect 28672 18650 28678 18737
rect 29024 18696 29070 18708
rect 29024 18650 29030 18696
rect 28672 18500 29030 18650
rect 28672 18252 28678 18500
rect 29024 18466 29030 18500
rect 29064 18650 29070 18696
rect 29540 18696 29586 18708
rect 29540 18650 29546 18696
rect 29064 18500 29546 18650
rect 29064 18466 29070 18500
rect 29024 18454 29070 18466
rect 29540 18466 29546 18500
rect 29580 18650 29586 18696
rect 30056 18696 30102 18708
rect 30056 18650 30062 18696
rect 29580 18500 30062 18650
rect 29580 18466 29586 18500
rect 29540 18454 29586 18466
rect 30056 18466 30062 18500
rect 30096 18650 30102 18696
rect 30572 18696 30618 18708
rect 30572 18650 30578 18696
rect 30096 18500 30578 18650
rect 30096 18466 30102 18500
rect 30056 18454 30102 18466
rect 30572 18466 30578 18500
rect 30612 18650 30618 18696
rect 31088 18696 31134 18708
rect 31088 18650 31094 18696
rect 30612 18500 31094 18650
rect 30612 18466 30618 18500
rect 30572 18454 30618 18466
rect 31088 18466 31094 18500
rect 31128 18650 31134 18696
rect 31604 18696 31650 18708
rect 31604 18650 31610 18696
rect 31128 18500 31610 18650
rect 31128 18466 31134 18500
rect 31088 18454 31134 18466
rect 31604 18466 31610 18500
rect 31644 18650 31650 18696
rect 32120 18696 32166 18708
rect 32120 18650 32126 18696
rect 31644 18500 32126 18650
rect 31644 18466 31650 18500
rect 31604 18454 31650 18466
rect 32120 18466 32126 18500
rect 32160 18650 32166 18696
rect 32160 18500 32170 18650
rect 32890 18538 32990 18760
rect 33850 18730 34730 18760
rect 33850 18710 34050 18730
rect 34300 18710 34730 18730
rect 32890 18504 32904 18538
rect 32972 18504 32990 18538
rect 32890 18500 32990 18504
rect 32160 18466 32166 18500
rect 32892 18498 32984 18500
rect 32120 18454 32166 18466
rect 33478 18492 33524 18504
rect 32836 18445 32882 18457
rect 28820 18390 32120 18410
rect 28820 18356 28834 18390
rect 29002 18356 29092 18390
rect 29260 18356 29350 18390
rect 29518 18356 29608 18390
rect 29776 18356 29866 18390
rect 30034 18356 30124 18390
rect 30292 18356 30382 18390
rect 30550 18356 30640 18390
rect 30808 18356 30898 18390
rect 31066 18356 31156 18390
rect 31324 18356 31414 18390
rect 31582 18356 31672 18390
rect 31840 18356 31930 18390
rect 32098 18356 32120 18390
rect 28820 18320 32120 18356
rect 32836 18330 32842 18445
rect 28480 18240 28678 18252
rect 28480 17990 28640 18240
rect 28480 17870 28500 17990
rect 28620 17870 28640 17990
rect 29670 18030 29760 18320
rect 32610 18315 32842 18330
rect 32610 18199 32708 18315
rect 32742 18199 32842 18315
rect 32610 18180 32842 18199
rect 29670 18020 32120 18030
rect 29670 17950 29680 18020
rect 29750 17998 32120 18020
rect 29750 17964 30124 17998
rect 30292 17964 30382 17998
rect 30550 17964 30640 17998
rect 30808 17964 30898 17998
rect 31066 17964 31156 17998
rect 31324 17964 31414 17998
rect 31582 17964 31672 17998
rect 31840 17964 31930 17998
rect 32098 17964 32120 17998
rect 29750 17950 32120 17964
rect 29670 17940 32120 17950
rect 28480 17570 28640 17870
rect 30056 17888 30102 17900
rect 30056 17658 30062 17888
rect 30096 17850 30102 17888
rect 30572 17888 30618 17900
rect 30572 17850 30578 17888
rect 30096 17700 30578 17850
rect 30096 17658 30102 17700
rect 30056 17646 30102 17658
rect 30572 17658 30578 17700
rect 30612 17850 30618 17888
rect 31088 17888 31134 17900
rect 31088 17850 31094 17888
rect 30612 17700 31094 17850
rect 30612 17658 30618 17700
rect 30572 17646 30618 17658
rect 31088 17658 31094 17700
rect 31128 17850 31134 17888
rect 31604 17888 31650 17900
rect 31604 17850 31610 17888
rect 31128 17700 31610 17850
rect 31128 17658 31134 17700
rect 31088 17646 31134 17658
rect 31604 17658 31610 17700
rect 31644 17850 31650 17888
rect 32120 17888 32166 17900
rect 32120 17850 32126 17888
rect 31644 17700 32126 17850
rect 31644 17658 31650 17700
rect 31604 17646 31650 17658
rect 32120 17658 32126 17700
rect 32160 17850 32166 17888
rect 32610 17850 32690 18180
rect 32836 18069 32842 18180
rect 32876 18069 32882 18445
rect 32836 18057 32882 18069
rect 32994 18445 33040 18457
rect 32994 18069 33000 18445
rect 33034 18330 33040 18445
rect 33478 18330 33484 18492
rect 33034 18310 33484 18330
rect 33034 18200 33230 18310
rect 33340 18200 33484 18310
rect 33034 18180 33484 18200
rect 33034 18069 33040 18180
rect 32994 18057 33040 18069
rect 33478 18079 33484 18180
rect 33518 18079 33524 18492
rect 33478 18067 33524 18079
rect 33636 18492 33682 18504
rect 33636 18079 33642 18492
rect 33676 18330 33682 18492
rect 33770 18400 33816 18412
rect 33770 18330 33776 18400
rect 33676 18180 33776 18330
rect 33676 18079 33682 18180
rect 33636 18067 33682 18079
rect 32892 18010 32984 18016
rect 32892 17976 32904 18010
rect 32972 17976 32984 18010
rect 32892 17970 32984 17976
rect 33530 18012 33630 18020
rect 33530 17978 33546 18012
rect 33614 17978 33630 18012
rect 32160 17700 32690 17850
rect 33530 17830 33630 17978
rect 33770 17874 33776 18180
rect 33810 18330 33816 18400
rect 33810 18310 34030 18330
rect 33810 18200 33890 18310
rect 34010 18200 34030 18310
rect 33810 18180 34030 18200
rect 33810 17874 33816 18180
rect 33870 17900 34030 18180
rect 34100 18310 34260 18330
rect 34100 18200 34120 18310
rect 34240 18200 34260 18310
rect 33770 17862 33816 17874
rect 33850 17880 34050 17900
rect 34100 17880 34260 18200
rect 34300 17880 34500 17900
rect 32160 17658 32166 17700
rect 32120 17646 32166 17658
rect 29922 17617 29968 17629
rect 28460 17540 28660 17570
rect 29922 17540 29928 17617
rect 28460 17390 29928 17540
rect 28460 17370 28660 17390
rect 28480 16720 28640 17370
rect 29922 17132 29928 17390
rect 29962 17540 29968 17617
rect 30314 17576 30360 17588
rect 30314 17540 30320 17576
rect 29962 17390 30320 17540
rect 29962 17132 29968 17390
rect 30314 17346 30320 17390
rect 30354 17540 30360 17576
rect 30830 17576 30876 17588
rect 30830 17540 30836 17576
rect 30354 17390 30836 17540
rect 30354 17346 30360 17390
rect 30314 17334 30360 17346
rect 30830 17346 30836 17390
rect 30870 17540 30876 17576
rect 31346 17576 31392 17588
rect 31346 17540 31352 17576
rect 30870 17390 31352 17540
rect 30870 17346 30876 17390
rect 30830 17334 30876 17346
rect 31346 17346 31352 17390
rect 31386 17540 31392 17576
rect 31862 17576 31908 17588
rect 31862 17540 31868 17576
rect 31386 17390 31868 17540
rect 31386 17346 31392 17390
rect 31346 17334 31392 17346
rect 31862 17346 31868 17390
rect 31902 17346 31908 17576
rect 31862 17334 31908 17346
rect 32610 17410 32690 17700
rect 33230 17770 33630 17830
rect 32892 17618 32984 17624
rect 32892 17584 32904 17618
rect 32972 17584 32984 17618
rect 32892 17578 32984 17584
rect 32836 17525 32882 17537
rect 32836 17410 32842 17525
rect 32610 17395 32842 17410
rect 32610 17279 32708 17395
rect 32742 17279 32842 17395
rect 30112 17270 30304 17276
rect 30112 17236 30124 17270
rect 30292 17236 30304 17270
rect 30112 17230 30304 17236
rect 30370 17270 30562 17276
rect 30370 17236 30382 17270
rect 30550 17236 30562 17270
rect 30370 17230 30562 17236
rect 30628 17270 30820 17276
rect 30628 17236 30640 17270
rect 30808 17236 30820 17270
rect 30628 17230 30820 17236
rect 30886 17270 31078 17276
rect 30886 17236 30898 17270
rect 31066 17236 31078 17270
rect 30886 17230 31078 17236
rect 31144 17270 31336 17276
rect 31144 17236 31156 17270
rect 31324 17236 31336 17270
rect 31144 17230 31336 17236
rect 31402 17270 31594 17276
rect 31402 17236 31414 17270
rect 31582 17236 31594 17270
rect 31402 17230 31594 17236
rect 31660 17270 31852 17276
rect 31660 17236 31672 17270
rect 31840 17236 31852 17270
rect 31660 17230 31852 17236
rect 31918 17270 32110 17276
rect 31918 17236 31930 17270
rect 32098 17236 32110 17270
rect 32610 17260 32842 17279
rect 31918 17230 32110 17236
rect 32836 17149 32842 17260
rect 32876 17149 32882 17525
rect 32836 17137 32882 17149
rect 32994 17525 33040 17537
rect 32994 17149 33000 17525
rect 33034 17410 33040 17525
rect 33230 17410 33330 17770
rect 33530 17622 33630 17770
rect 33530 17588 33546 17622
rect 33614 17588 33630 17622
rect 33530 17580 33630 17588
rect 33770 17726 33816 17738
rect 33478 17521 33524 17533
rect 33478 17410 33484 17521
rect 33034 17260 33484 17410
rect 33034 17149 33040 17260
rect 32994 17137 33040 17149
rect 29922 17120 29968 17132
rect 33478 17108 33484 17260
rect 33518 17108 33524 17521
rect 32890 17090 32990 17100
rect 33478 17096 33524 17108
rect 33636 17521 33682 17533
rect 33636 17108 33642 17521
rect 33676 17410 33682 17521
rect 33770 17410 33776 17726
rect 33676 17260 33776 17410
rect 33676 17108 33682 17260
rect 33770 17200 33776 17260
rect 33810 17410 33816 17726
rect 33850 17720 34500 17880
rect 33850 17700 34050 17720
rect 34300 17700 34500 17720
rect 33870 17410 34030 17700
rect 33810 17260 34030 17410
rect 33810 17200 33816 17260
rect 33770 17188 33816 17200
rect 33636 17096 33682 17108
rect 32890 17056 32904 17090
rect 32972 17056 32990 17090
rect 29922 16972 29968 16984
rect 29922 16720 29928 16972
rect 28480 16570 29928 16720
rect 29922 16487 29928 16570
rect 29962 16720 29968 16972
rect 30112 16868 30304 16874
rect 30112 16834 30124 16868
rect 30292 16834 30304 16868
rect 30112 16828 30304 16834
rect 30370 16868 30562 16874
rect 30370 16834 30382 16868
rect 30550 16834 30562 16868
rect 30370 16828 30562 16834
rect 30628 16868 30820 16874
rect 30628 16834 30640 16868
rect 30808 16834 30820 16868
rect 30628 16828 30820 16834
rect 30886 16868 31078 16874
rect 30886 16834 30898 16868
rect 31066 16834 31078 16868
rect 30886 16828 31078 16834
rect 31144 16868 31336 16874
rect 31144 16834 31156 16868
rect 31324 16834 31336 16868
rect 31144 16828 31336 16834
rect 31402 16868 31594 16874
rect 31402 16834 31414 16868
rect 31582 16834 31594 16868
rect 31402 16828 31594 16834
rect 31660 16868 31852 16874
rect 31660 16834 31672 16868
rect 31840 16834 31852 16868
rect 31660 16828 31852 16834
rect 31918 16868 32110 16874
rect 31918 16834 31930 16868
rect 32098 16834 32110 16868
rect 31918 16828 32110 16834
rect 32890 16840 32990 17056
rect 33870 17020 34030 17040
rect 33870 16910 33890 17020
rect 34010 16910 34030 17020
rect 33870 16890 34030 16910
rect 33850 16840 34050 16890
rect 30056 16758 30102 16770
rect 30056 16720 30062 16758
rect 29962 16570 30062 16720
rect 29962 16487 29968 16570
rect 30056 16528 30062 16570
rect 30096 16720 30102 16758
rect 30572 16758 30618 16770
rect 30572 16720 30578 16758
rect 30096 16570 30578 16720
rect 30096 16528 30102 16570
rect 30056 16516 30102 16528
rect 30572 16528 30578 16570
rect 30612 16720 30618 16758
rect 31088 16758 31134 16770
rect 31088 16720 31094 16758
rect 30612 16570 31094 16720
rect 30612 16528 30618 16570
rect 30572 16516 30618 16528
rect 31088 16528 31094 16570
rect 31128 16720 31134 16758
rect 31604 16758 31650 16770
rect 31604 16720 31610 16758
rect 31128 16570 31610 16720
rect 31128 16528 31134 16570
rect 31088 16516 31134 16528
rect 31604 16528 31610 16570
rect 31644 16720 31650 16758
rect 32120 16758 32166 16770
rect 32120 16720 32126 16758
rect 31644 16570 32126 16720
rect 31644 16528 31650 16570
rect 31604 16516 31650 16528
rect 32120 16528 32126 16570
rect 32160 16528 32166 16758
rect 32890 16740 34050 16840
rect 33850 16690 34050 16740
rect 32120 16516 32166 16528
rect 29922 16475 29968 16487
rect 30314 16446 30360 16458
rect 28460 16410 28660 16440
rect 30314 16410 30320 16446
rect 28460 16380 30320 16410
rect 28460 16290 29670 16380
rect 29760 16290 30320 16380
rect 28460 16260 30320 16290
rect 28460 16240 28660 16260
rect 28480 15990 28640 16240
rect 29670 16170 29760 16260
rect 30314 16216 30320 16260
rect 30354 16410 30360 16446
rect 30830 16446 30876 16458
rect 30830 16410 30836 16446
rect 30354 16260 30836 16410
rect 30354 16216 30360 16260
rect 30314 16204 30360 16216
rect 30830 16216 30836 16260
rect 30870 16410 30876 16446
rect 31346 16446 31392 16458
rect 31346 16410 31352 16446
rect 30870 16260 31352 16410
rect 30870 16216 30876 16260
rect 30830 16204 30876 16216
rect 31346 16216 31352 16260
rect 31386 16410 31392 16446
rect 31862 16446 31908 16458
rect 31862 16410 31868 16446
rect 31386 16260 31868 16410
rect 31386 16216 31392 16260
rect 31346 16204 31392 16216
rect 31862 16216 31868 16260
rect 31902 16410 31908 16446
rect 31902 16260 31910 16410
rect 31902 16216 31908 16260
rect 31862 16204 31908 16216
rect 29670 16140 32120 16170
rect 29670 16106 30124 16140
rect 30292 16106 30382 16140
rect 30550 16106 30640 16140
rect 30808 16106 30898 16140
rect 31066 16106 31156 16140
rect 31324 16106 31414 16140
rect 31582 16106 31672 16140
rect 31840 16106 31930 16140
rect 32098 16106 32120 16140
rect 29670 16080 32120 16106
rect 33534 16112 33626 16118
rect 33534 16078 33546 16112
rect 33614 16078 33626 16112
rect 33534 16072 33626 16078
rect 28460 15790 28660 15990
rect 28480 15530 28640 15790
rect 34530 15530 34730 15550
rect 28480 15370 34730 15530
rect 34530 15350 34730 15370
<< via1 >>
rect 1040 32980 1160 33100
rect 10180 32980 10300 33100
rect 19370 32980 19490 33100
rect 1600 25940 1720 26060
rect 4120 26060 4280 26220
rect 9660 26080 9780 26180
rect 3520 22700 3680 22860
rect 10740 25940 10860 26060
rect 13260 26060 13420 26220
rect 18800 26080 18920 26180
rect 12660 22700 12820 22860
rect 19930 25940 20050 26060
rect 22450 26060 22610 26220
rect 27990 26080 28110 26180
rect 33890 26080 34010 26200
rect 32380 25320 32470 25410
rect 28500 23030 28620 23150
rect 21850 22700 22010 22860
rect 12660 22080 12810 22240
rect 21830 22080 22010 22240
rect 28720 22080 28870 22240
rect 33690 20050 33790 20160
rect 33890 19740 34010 19850
rect 32800 19540 32890 19630
rect 28500 17870 28620 17990
rect 29680 17950 29750 18020
rect 33230 18200 33340 18310
rect 33890 18200 34010 18310
rect 34120 18200 34240 18310
rect 33890 16910 34010 17020
rect 29670 16290 29760 16380
<< metal2 >>
rect 1040 33100 1160 33110
rect 1040 32970 1160 32980
rect 10180 33100 10300 33110
rect 10180 32970 10300 32980
rect 19370 33100 19490 33110
rect 19370 32970 19490 32980
rect 4120 26220 4280 26230
rect 1600 26060 1720 26070
rect 13260 26220 13420 26230
rect 9660 26180 9780 26190
rect 9660 26070 9780 26080
rect 4120 26050 4280 26060
rect 10740 26060 10860 26070
rect 1600 25930 1720 25940
rect 22450 26220 22610 26230
rect 18800 26180 18920 26190
rect 18800 26070 18920 26080
rect 13260 26050 13420 26060
rect 19930 26060 20050 26070
rect 10740 25930 10860 25940
rect 33890 26200 34010 26210
rect 27990 26180 28110 26190
rect 27990 26070 28110 26080
rect 33890 26070 34010 26080
rect 22450 26050 22610 26060
rect 19930 25930 20050 25940
rect 32490 25420 34260 25430
rect 32360 25410 34260 25420
rect 32360 25320 32380 25410
rect 32470 25320 34260 25410
rect 32360 25300 34260 25320
rect 28480 23150 28640 23170
rect 28480 23030 28500 23150
rect 28620 23030 28640 23150
rect 3520 22860 3680 22870
rect 3520 22690 3680 22700
rect 12660 22860 12820 22870
rect 12660 22690 12820 22700
rect 21850 22860 22010 22870
rect 21850 22690 22010 22700
rect 12640 22240 22030 22260
rect 12640 22080 12660 22240
rect 12810 22080 21830 22240
rect 22010 22080 22030 22240
rect 12640 22060 22030 22080
rect 28480 17990 28640 23030
rect 34100 22260 34260 25300
rect 28700 22240 34260 22260
rect 28700 22080 28720 22240
rect 28870 22080 34260 22240
rect 28700 22060 34260 22080
rect 33690 20160 33790 20170
rect 33690 20040 33790 20050
rect 33870 19850 34030 19870
rect 33870 19740 33890 19850
rect 34010 19740 34030 19850
rect 32790 19630 32900 19640
rect 32790 19540 32800 19630
rect 32890 19540 32900 19630
rect 32790 19020 32900 19540
rect 32790 18910 33340 19020
rect 33230 18310 33340 18910
rect 33230 18190 33340 18200
rect 33870 18310 34030 19740
rect 33870 18200 33890 18310
rect 34010 18200 34030 18310
rect 33870 18180 34030 18200
rect 34100 18310 34260 22060
rect 34100 18200 34120 18310
rect 34240 18200 34260 18310
rect 34100 18180 34260 18200
rect 28480 17870 28500 17990
rect 28620 17870 28640 17990
rect 28480 17860 28640 17870
rect 29670 18020 29760 18030
rect 29670 17950 29680 18020
rect 29750 17950 29760 18020
rect 29670 16380 29760 17950
rect 33890 17020 34010 17030
rect 33890 16900 34010 16910
rect 29670 16280 29760 16290
<< via2 >>
rect 1040 32980 1160 33100
rect 10180 32980 10300 33100
rect 19370 32980 19490 33100
rect 1600 25940 1720 26060
rect 4120 26060 4280 26220
rect 9660 26080 9780 26180
rect 10740 25940 10860 26060
rect 13260 26060 13420 26220
rect 18800 26080 18920 26180
rect 19930 25940 20050 26060
rect 22450 26060 22610 26220
rect 27990 26080 28110 26180
rect 33890 26080 34010 26200
rect 3520 22700 3680 22860
rect 12660 22700 12820 22860
rect 21850 22700 22010 22860
rect 33690 20050 33790 20160
rect 32800 19540 32890 19630
rect 33890 16910 34010 17020
<< metal3 >>
rect 1030 33100 1170 33105
rect 1030 32980 1040 33100
rect 1160 32980 1170 33100
rect 1030 32975 1170 32980
rect 10170 33100 10310 33105
rect 10170 32980 10180 33100
rect 10300 32980 10310 33100
rect 10170 32975 10310 32980
rect 19360 33100 19500 33105
rect 19360 32980 19370 33100
rect 19490 32980 19500 33100
rect 19360 32975 19500 32980
rect 1100 32752 7399 32780
rect 1100 26608 1120 32752
rect 1184 26608 7399 32752
rect 1100 26580 7399 26608
rect 10240 32752 16539 32780
rect 10240 26608 10260 32752
rect 10324 26608 16539 32752
rect 10240 26580 16539 26608
rect 19430 32752 25729 32780
rect 19430 26608 19450 32752
rect 19514 26608 25729 32752
rect 19430 26580 25729 26608
rect 4110 26220 4290 26225
rect 1590 26060 1730 26065
rect 1590 25940 1600 26060
rect 1720 25940 1730 26060
rect 4110 26060 4120 26220
rect 4280 26060 4290 26220
rect 13250 26220 13430 26225
rect 9650 26180 9790 26185
rect 9650 26080 9660 26180
rect 9780 26080 9790 26180
rect 9650 26075 9790 26080
rect 4110 26055 4290 26060
rect 10730 26060 10870 26065
rect 1590 25935 1730 25940
rect 3700 25922 9999 25950
rect 10730 25940 10740 26060
rect 10860 25940 10870 26060
rect 13250 26060 13260 26220
rect 13420 26060 13430 26220
rect 22440 26220 22620 26225
rect 18790 26180 18930 26185
rect 18790 26080 18800 26180
rect 18920 26080 18930 26180
rect 18790 26075 18930 26080
rect 13250 26055 13430 26060
rect 19920 26060 20060 26065
rect 10730 25935 10870 25940
rect 3700 22885 3720 25922
rect 3690 22865 3720 22885
rect 3510 22860 3720 22865
rect 3510 22700 3520 22860
rect 3680 22700 3720 22860
rect 3510 22695 3720 22700
rect 3690 22675 3720 22695
rect 3700 19778 3720 22675
rect 3784 19778 9999 25922
rect 12840 25922 19139 25950
rect 19920 25940 19930 26060
rect 20050 25940 20060 26060
rect 22440 26060 22450 26220
rect 22610 26060 22620 26220
rect 33870 26200 34030 26220
rect 27980 26180 28120 26185
rect 27980 26080 27990 26180
rect 28110 26080 28120 26180
rect 27980 26075 28120 26080
rect 33870 26080 33890 26200
rect 34010 26080 34030 26200
rect 22440 26055 22620 26060
rect 19920 25935 20060 25940
rect 12840 22885 12860 25922
rect 12830 22865 12860 22885
rect 12650 22860 12860 22865
rect 12650 22700 12660 22860
rect 12820 22700 12860 22860
rect 12650 22695 12860 22700
rect 12830 22675 12860 22695
rect 3700 19750 9999 19778
rect 12840 19778 12860 22675
rect 12924 19778 19139 25922
rect 22030 25922 28329 25950
rect 22030 22885 22050 25922
rect 22020 22865 22050 22885
rect 21840 22860 22050 22865
rect 21840 22700 21850 22860
rect 22010 22700 22050 22860
rect 21840 22695 22050 22700
rect 22020 22675 22050 22695
rect 12840 19750 19139 19778
rect 22030 19778 22050 22675
rect 22114 19778 28329 25922
rect 28890 25302 33789 25330
rect 28890 20558 33705 25302
rect 33769 20558 33789 25302
rect 28890 20530 33789 20558
rect 33680 20160 33800 20165
rect 33680 20050 33690 20160
rect 33790 20050 33800 20160
rect 33680 20045 33800 20050
rect 22030 19750 28329 19778
rect 3700 19622 9999 19650
rect 3700 13478 3720 19622
rect 3784 13478 9999 19622
rect 3700 13450 9999 13478
rect 12840 19622 19139 19650
rect 12840 13478 12860 19622
rect 12924 13478 19139 19622
rect 12840 13450 19139 13478
rect 22030 19622 28329 19650
rect 22030 13478 22050 19622
rect 22114 13478 28329 19622
rect 32790 19630 32900 19635
rect 32790 19540 32800 19630
rect 32890 19540 32900 19630
rect 32790 19535 32900 19540
rect 33870 17020 34030 26080
rect 33870 16910 33890 17020
rect 34010 16910 34030 17020
rect 33870 16890 34030 16910
rect 22030 13450 28329 13478
rect 3700 13322 9999 13350
rect 3700 7178 3720 13322
rect 3784 7178 9999 13322
rect 3700 7150 9999 7178
rect 12840 13322 19139 13350
rect 12840 7178 12860 13322
rect 12924 7178 19139 13322
rect 12840 7150 19139 7178
rect 22030 13322 28329 13350
rect 22030 7178 22050 13322
rect 22114 7178 28329 13322
rect 22030 7150 28329 7178
<< via3 >>
rect 1040 32980 1160 33100
rect 10180 32980 10300 33100
rect 19370 32980 19490 33100
rect 1120 26608 1184 32752
rect 10260 26608 10324 32752
rect 19450 26608 19514 32752
rect 1600 25940 1720 26060
rect 4120 26060 4280 26220
rect 9660 26080 9780 26180
rect 10740 25940 10860 26060
rect 13260 26060 13420 26220
rect 18800 26080 18920 26180
rect 3520 22700 3680 22860
rect 3720 19778 3784 25922
rect 19930 25940 20050 26060
rect 22450 26060 22610 26220
rect 27990 26080 28110 26180
rect 12660 22700 12820 22860
rect 12860 19778 12924 25922
rect 21850 22700 22010 22860
rect 22050 19778 22114 25922
rect 33705 20558 33769 25302
rect 33690 20050 33790 20160
rect 3720 13478 3784 19622
rect 12860 13478 12924 19622
rect 22050 13478 22114 19622
rect 32800 19540 32890 19630
rect 3720 7178 3784 13322
rect 12860 7178 12924 13322
rect 22050 7178 22114 13322
<< mimcap >>
rect 1299 32640 7299 32680
rect 1299 26720 1339 32640
rect 7259 26720 7299 32640
rect 1299 26680 7299 26720
rect 10439 32640 16439 32680
rect 10439 26720 10479 32640
rect 16399 26720 16439 32640
rect 10439 26680 16439 26720
rect 19629 32640 25629 32680
rect 19629 26720 19669 32640
rect 25589 26720 25629 32640
rect 19629 26680 25629 26720
rect 3899 25810 9899 25850
rect 3899 19890 3939 25810
rect 9859 19890 9899 25810
rect 3899 19850 9899 19890
rect 13039 25810 19039 25850
rect 13039 19890 13079 25810
rect 18999 19890 19039 25810
rect 13039 19850 19039 19890
rect 22229 25810 28229 25850
rect 22229 19890 22269 25810
rect 28189 19890 28229 25810
rect 28990 25190 33590 25230
rect 28990 20670 29030 25190
rect 33550 20670 33590 25190
rect 28990 20630 33590 20670
rect 22229 19850 28229 19890
rect 3899 19510 9899 19550
rect 3899 13590 3939 19510
rect 9859 13590 9899 19510
rect 3899 13550 9899 13590
rect 13039 19510 19039 19550
rect 13039 13590 13079 19510
rect 18999 13590 19039 19510
rect 13039 13550 19039 13590
rect 22229 19510 28229 19550
rect 22229 13590 22269 19510
rect 28189 13590 28229 19510
rect 22229 13550 28229 13590
rect 3899 13210 9899 13250
rect 3899 7290 3939 13210
rect 9859 7290 9899 13210
rect 3899 7250 9899 7290
rect 13039 13210 19039 13250
rect 13039 7290 13079 13210
rect 18999 7290 19039 13210
rect 13039 7250 19039 7290
rect 22229 13210 28229 13250
rect 22229 7290 22269 13210
rect 28189 7290 28229 13210
rect 22229 7250 28229 7290
<< mimcapcontact >>
rect 1339 26720 7259 32640
rect 10479 26720 16399 32640
rect 19669 26720 25589 32640
rect 3939 19890 9859 25810
rect 13079 19890 18999 25810
rect 22269 19890 28189 25810
rect 29030 20670 33550 25190
rect 3939 13590 9859 19510
rect 13079 13590 18999 19510
rect 22269 13590 28189 19510
rect 3939 7290 9859 13210
rect 13079 7290 18999 13210
rect 22269 7290 28189 13210
<< metal4 >>
rect 1039 33100 1161 33101
rect 1039 32980 1040 33100
rect 1160 32980 1161 33100
rect 1039 32979 1161 32980
rect 10179 33100 10301 33101
rect 10179 32980 10180 33100
rect 10300 32980 10301 33100
rect 10179 32979 10301 32980
rect 19369 33100 19491 33101
rect 19369 32980 19370 33100
rect 19490 32980 19491 33100
rect 19369 32979 19491 32980
rect 1060 32880 1160 32979
rect 10200 32880 10300 32979
rect 19390 32880 19490 32979
rect 1060 32780 1200 32880
rect 10200 32780 10340 32880
rect 19390 32780 19530 32880
rect 1100 32752 1200 32780
rect 1100 32720 1120 32752
rect 1104 26608 1120 32720
rect 1184 26608 1200 32752
rect 10240 32752 10340 32780
rect 10240 32720 10260 32752
rect 1338 32640 7260 32641
rect 1338 26720 1339 32640
rect 7259 26720 7260 32640
rect 1338 26719 7260 26720
rect 1104 26592 1200 26608
rect 1580 26060 1740 26719
rect 10244 26608 10260 32720
rect 10324 26608 10340 32752
rect 19430 32752 19530 32780
rect 19430 32720 19450 32752
rect 10478 32640 16400 32641
rect 10478 26720 10479 32640
rect 16399 26720 16400 32640
rect 10478 26719 16400 26720
rect 10244 26592 10340 26608
rect 1580 25940 1600 26060
rect 1720 25940 1740 26060
rect 4100 26220 4300 26240
rect 4100 26060 4120 26220
rect 4280 26060 4300 26220
rect 1580 25920 1740 25940
rect 3727 25938 3831 26000
rect 3704 25922 3831 25938
rect 3704 22880 3720 25922
rect 3500 22860 3720 22880
rect 3500 22700 3520 22860
rect 3680 22700 3720 22860
rect 3500 22680 3720 22700
rect 3704 19778 3720 22680
rect 3784 19778 3831 25922
rect 4100 25811 4300 26060
rect 9640 26180 9800 26200
rect 9640 26080 9660 26180
rect 9780 26080 9800 26180
rect 6847 25811 6951 26000
rect 9640 25811 9800 26080
rect 10720 26060 10880 26719
rect 19434 26608 19450 32720
rect 19514 26608 19530 32752
rect 19668 32640 25590 32641
rect 19668 26720 19669 32640
rect 25589 26720 25590 32640
rect 19668 26719 25590 26720
rect 19434 26592 19530 26608
rect 10720 25940 10740 26060
rect 10860 25940 10880 26060
rect 13240 26220 13440 26240
rect 13240 26060 13260 26220
rect 13420 26060 13440 26220
rect 10720 25920 10880 25940
rect 12867 25938 12971 26000
rect 12844 25922 12971 25938
rect 3938 25810 9860 25811
rect 3938 19890 3939 25810
rect 9859 19890 9860 25810
rect 12844 22880 12860 25922
rect 12640 22860 12860 22880
rect 12640 22700 12660 22860
rect 12820 22700 12860 22860
rect 12640 22680 12860 22700
rect 3938 19889 9860 19890
rect 3704 19762 3831 19778
rect 3727 19638 3831 19762
rect 3704 19622 3831 19638
rect 3704 13478 3720 19622
rect 3784 13478 3831 19622
rect 6847 19511 6951 19889
rect 12844 19778 12860 22680
rect 12924 19778 12971 25922
rect 13240 25811 13440 26060
rect 18780 26180 18940 26200
rect 18780 26080 18800 26180
rect 18920 26080 18940 26180
rect 15987 25811 16091 26000
rect 18780 25811 18940 26080
rect 19910 26060 20070 26719
rect 19910 25940 19930 26060
rect 20050 25940 20070 26060
rect 22430 26220 22630 26240
rect 22430 26060 22450 26220
rect 22610 26060 22630 26220
rect 19910 25920 20070 25940
rect 22057 25938 22161 26000
rect 22034 25922 22161 25938
rect 13078 25810 19000 25811
rect 13078 19890 13079 25810
rect 18999 19890 19000 25810
rect 22034 22880 22050 25922
rect 21830 22860 22050 22880
rect 21830 22700 21850 22860
rect 22010 22700 22050 22860
rect 21830 22680 22050 22700
rect 13078 19889 19000 19890
rect 12844 19762 12971 19778
rect 12867 19638 12971 19762
rect 12844 19622 12971 19638
rect 3938 19510 9860 19511
rect 3938 13590 3939 19510
rect 9859 13590 9860 19510
rect 3938 13589 9860 13590
rect 3704 13462 3831 13478
rect 3727 13338 3831 13462
rect 3704 13322 3831 13338
rect 3704 7178 3720 13322
rect 3784 7178 3831 13322
rect 6847 13211 6951 13589
rect 12844 13478 12860 19622
rect 12924 13478 12971 19622
rect 15987 19511 16091 19889
rect 22034 19778 22050 22680
rect 22114 19778 22161 25922
rect 22430 25811 22630 26060
rect 27970 26180 28130 26200
rect 27970 26080 27990 26180
rect 28110 26080 28130 26180
rect 25177 25811 25281 26000
rect 27970 25811 28130 26080
rect 22268 25810 28190 25811
rect 22268 19890 22269 25810
rect 28189 19890 28190 25810
rect 33689 25302 33785 25318
rect 29029 25190 33551 25191
rect 29029 20670 29030 25190
rect 33550 20670 33551 25190
rect 29029 20669 33551 20670
rect 22268 19889 28190 19890
rect 22034 19762 22161 19778
rect 22057 19638 22161 19762
rect 22034 19622 22161 19638
rect 13078 19510 19000 19511
rect 13078 13590 13079 19510
rect 18999 13590 19000 19510
rect 13078 13589 19000 13590
rect 12844 13462 12971 13478
rect 12867 13338 12971 13462
rect 12844 13322 12971 13338
rect 3938 13210 9860 13211
rect 3938 7290 3939 13210
rect 9859 7290 9860 13210
rect 3938 7289 9860 7290
rect 3704 7162 3831 7178
rect 3727 7100 3831 7162
rect 6847 7100 6951 7289
rect 12844 7178 12860 13322
rect 12924 7178 12971 13322
rect 15987 13211 16091 13589
rect 22034 13478 22050 19622
rect 22114 13478 22161 19622
rect 25177 19511 25281 19889
rect 32790 19630 32900 20669
rect 33689 20558 33705 25302
rect 33769 20570 33785 25302
rect 33769 20558 33790 20570
rect 33689 20542 33790 20558
rect 33690 20161 33790 20542
rect 33689 20160 33791 20161
rect 33689 20050 33690 20160
rect 33790 20050 33791 20160
rect 33689 20049 33791 20050
rect 32790 19540 32800 19630
rect 32890 19540 32900 19630
rect 32790 19530 32900 19540
rect 22268 19510 28190 19511
rect 22268 13590 22269 19510
rect 28189 13590 28190 19510
rect 22268 13589 28190 13590
rect 22034 13462 22161 13478
rect 22057 13338 22161 13462
rect 22034 13322 22161 13338
rect 13078 13210 19000 13211
rect 13078 7290 13079 13210
rect 18999 7290 19000 13210
rect 13078 7289 19000 7290
rect 12844 7162 12971 7178
rect 12867 7100 12971 7162
rect 15987 7100 16091 7289
rect 22034 7178 22050 13322
rect 22114 7178 22161 13322
rect 25177 13211 25281 13589
rect 22268 13210 28190 13211
rect 22268 7290 22269 13210
rect 28189 7290 28190 13210
rect 22268 7289 28190 7290
rect 22034 7162 22161 7178
rect 22057 7100 22161 7162
rect 25177 7100 25281 7289
<< labels >>
flabel metal1 770 33120 970 33320 0 FreeSans 256 0 0 0 top_in
port 0 nsew
flabel metal1 770 22680 970 22880 0 FreeSans 256 0 0 0 top_gnd
port 1 nsew
flabel metal1 34530 15350 34730 15550 0 FreeSans 256 0 0 0 top_ibias
port 2 nsew
flabel metal1 34530 18710 34730 18910 0 FreeSans 256 0 0 0 top_ref
port 3 nsew
flabel metal1 34560 26040 34760 26240 0 FreeSans 256 0 0 0 top_out
port 4 nsew
flabel metal1 28460 15790 28660 15990 0 FreeSans 256 0 0 0 x4.ldo_ibias
flabel metal1 28460 26040 28660 26240 0 FreeSans 256 0 0 0 x4.ldo_in
flabel metal1 34300 18710 34500 18910 0 FreeSans 256 0 0 0 x4.ldo_ref
flabel metal1 34300 17700 34500 17900 0 FreeSans 256 0 0 0 x4.ldo_gnd
flabel metal1 34330 26040 34530 26240 0 FreeSans 256 0 0 0 x4.ldo_out
flabel metal1 28460 17370 28660 17570 0 FreeSans 256 0 0 0 x4.x1.VDD
flabel metal1 28460 16240 28660 16440 0 FreeSans 256 0 0 0 x4.x1.Ibias
flabel metal1 33850 17700 34050 17900 0 FreeSans 256 0 0 0 x4.x1.VSS
flabel metal1 33850 20010 34050 20210 0 FreeSans 256 0 0 0 x4.x1.Vout
flabel metal1 33850 18710 34050 18910 0 FreeSans 256 0 0 0 x4.x1.Vip
flabel metal1 33850 16690 34050 16890 0 FreeSans 256 0 0 0 x4.x1.Vin
flabel metal1 19330 22680 19530 22880 0 FreeSans 256 0 0 0 x3.ground
flabel metal1 19330 33120 19530 33320 0 FreeSans 256 0 0 0 x3.i
flabel metal1 28230 26040 28430 26240 0 FreeSans 256 0 0 0 x3.o
flabel metal1 10140 22680 10340 22880 0 FreeSans 256 0 0 0 x2.ground
flabel metal1 10140 33120 10340 33320 0 FreeSans 256 0 0 0 x2.i
flabel metal1 19040 26040 19240 26240 0 FreeSans 256 0 0 0 x2.o
flabel metal1 1000 22680 1200 22880 0 FreeSans 256 0 0 0 x1.ground
flabel metal1 1000 33120 1200 33320 0 FreeSans 256 0 0 0 x1.i
flabel metal1 9900 26040 10100 26240 0 FreeSans 256 0 0 0 x1.o
<< end >>
