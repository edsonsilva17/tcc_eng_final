magic
tech sky130A
timestamp 1712847951
<< pwell >>
rect -551 -279 551 279
<< mvnmos >>
rect -437 -150 -337 150
rect -308 -150 -208 150
rect -179 -150 -79 150
rect -50 -150 50 150
rect 79 -150 179 150
rect 208 -150 308 150
rect 337 -150 437 150
<< mvndiff >>
rect -466 144 -437 150
rect -466 -144 -460 144
rect -443 -144 -437 144
rect -466 -150 -437 -144
rect -337 144 -308 150
rect -337 -144 -331 144
rect -314 -144 -308 144
rect -337 -150 -308 -144
rect -208 144 -179 150
rect -208 -144 -202 144
rect -185 -144 -179 144
rect -208 -150 -179 -144
rect -79 144 -50 150
rect -79 -144 -73 144
rect -56 -144 -50 144
rect -79 -150 -50 -144
rect 50 144 79 150
rect 50 -144 56 144
rect 73 -144 79 144
rect 50 -150 79 -144
rect 179 144 208 150
rect 179 -144 185 144
rect 202 -144 208 144
rect 179 -150 208 -144
rect 308 144 337 150
rect 308 -144 314 144
rect 331 -144 337 144
rect 308 -150 337 -144
rect 437 144 466 150
rect 437 -144 443 144
rect 460 -144 466 144
rect 437 -150 466 -144
<< mvndiffc >>
rect -460 -144 -443 144
rect -331 -144 -314 144
rect -202 -144 -185 144
rect -73 -144 -56 144
rect 56 -144 73 144
rect 185 -144 202 144
rect 314 -144 331 144
rect 443 -144 460 144
<< mvpsubdiff >>
rect -533 255 533 261
rect -533 238 -479 255
rect 479 238 533 255
rect -533 232 533 238
rect -533 207 -504 232
rect -533 -207 -527 207
rect -510 -207 -504 207
rect 504 207 533 232
rect -533 -232 -504 -207
rect 504 -207 510 207
rect 527 -207 533 207
rect 504 -232 533 -207
rect -533 -238 533 -232
rect -533 -255 -479 -238
rect 479 -255 533 -238
rect -533 -261 533 -255
<< mvpsubdiffcont >>
rect -479 238 479 255
rect -527 -207 -510 207
rect 510 -207 527 207
rect -479 -255 479 -238
<< poly >>
rect -437 186 -337 194
rect -437 169 -429 186
rect -345 169 -337 186
rect -437 150 -337 169
rect -308 186 -208 194
rect -308 169 -300 186
rect -216 169 -208 186
rect -308 150 -208 169
rect -179 186 -79 194
rect -179 169 -171 186
rect -87 169 -79 186
rect -179 150 -79 169
rect -50 186 50 194
rect -50 169 -42 186
rect 42 169 50 186
rect -50 150 50 169
rect 79 186 179 194
rect 79 169 87 186
rect 171 169 179 186
rect 79 150 179 169
rect 208 186 308 194
rect 208 169 216 186
rect 300 169 308 186
rect 208 150 308 169
rect 337 186 437 194
rect 337 169 345 186
rect 429 169 437 186
rect 337 150 437 169
rect -437 -169 -337 -150
rect -437 -186 -429 -169
rect -345 -186 -337 -169
rect -437 -194 -337 -186
rect -308 -169 -208 -150
rect -308 -186 -300 -169
rect -216 -186 -208 -169
rect -308 -194 -208 -186
rect -179 -169 -79 -150
rect -179 -186 -171 -169
rect -87 -186 -79 -169
rect -179 -194 -79 -186
rect -50 -169 50 -150
rect -50 -186 -42 -169
rect 42 -186 50 -169
rect -50 -194 50 -186
rect 79 -169 179 -150
rect 79 -186 87 -169
rect 171 -186 179 -169
rect 79 -194 179 -186
rect 208 -169 308 -150
rect 208 -186 216 -169
rect 300 -186 308 -169
rect 208 -194 308 -186
rect 337 -169 437 -150
rect 337 -186 345 -169
rect 429 -186 437 -169
rect 337 -194 437 -186
<< polycont >>
rect -429 169 -345 186
rect -300 169 -216 186
rect -171 169 -87 186
rect -42 169 42 186
rect 87 169 171 186
rect 216 169 300 186
rect 345 169 429 186
rect -429 -186 -345 -169
rect -300 -186 -216 -169
rect -171 -186 -87 -169
rect -42 -186 42 -169
rect 87 -186 171 -169
rect 216 -186 300 -169
rect 345 -186 429 -169
<< locali >>
rect -527 238 -479 255
rect 479 238 527 255
rect -527 207 -510 238
rect 510 207 527 238
rect -437 169 -429 186
rect -345 169 -337 186
rect -308 169 -300 186
rect -216 169 -208 186
rect -179 169 -171 186
rect -87 169 -79 186
rect -50 169 -42 186
rect 42 169 50 186
rect 79 169 87 186
rect 171 169 179 186
rect 208 169 216 186
rect 300 169 308 186
rect 337 169 345 186
rect 429 169 437 186
rect -460 144 -443 152
rect -460 -152 -443 -144
rect -331 144 -314 152
rect -331 -152 -314 -144
rect -202 144 -185 152
rect -202 -152 -185 -144
rect -73 144 -56 152
rect -73 -152 -56 -144
rect 56 144 73 152
rect 56 -152 73 -144
rect 185 144 202 152
rect 185 -152 202 -144
rect 314 144 331 152
rect 314 -152 331 -144
rect 443 144 460 152
rect 443 -152 460 -144
rect -437 -186 -429 -169
rect -345 -186 -337 -169
rect -308 -186 -300 -169
rect -216 -186 -208 -169
rect -179 -186 -171 -169
rect -87 -186 -79 -169
rect -50 -186 -42 -169
rect 42 -186 50 -169
rect 79 -186 87 -169
rect 171 -186 179 -169
rect 208 -186 216 -169
rect 300 -186 308 -169
rect 337 -186 345 -169
rect 429 -186 437 -169
rect -527 -238 -510 -207
rect 510 -238 527 -207
rect -527 -255 -479 -238
rect 479 -255 527 -238
<< viali >>
rect -429 169 -345 186
rect -300 169 -216 186
rect -171 169 -87 186
rect -42 169 42 186
rect 87 169 171 186
rect 216 169 300 186
rect 345 169 429 186
rect -460 -144 -443 144
rect -331 -144 -314 144
rect -202 -144 -185 144
rect -73 -144 -56 144
rect 56 -144 73 144
rect 185 -144 202 144
rect 314 -144 331 144
rect 443 -144 460 144
rect -429 -186 -345 -169
rect -300 -186 -216 -169
rect -171 -186 -87 -169
rect -42 -186 42 -169
rect 87 -186 171 -169
rect 216 -186 300 -169
rect 345 -186 429 -169
<< metal1 >>
rect -435 186 -339 189
rect -435 169 -429 186
rect -345 169 -339 186
rect -435 166 -339 169
rect -306 186 -210 189
rect -306 169 -300 186
rect -216 169 -210 186
rect -306 166 -210 169
rect -177 186 -81 189
rect -177 169 -171 186
rect -87 169 -81 186
rect -177 166 -81 169
rect -48 186 48 189
rect -48 169 -42 186
rect 42 169 48 186
rect -48 166 48 169
rect 81 186 177 189
rect 81 169 87 186
rect 171 169 177 186
rect 81 166 177 169
rect 210 186 306 189
rect 210 169 216 186
rect 300 169 306 186
rect 210 166 306 169
rect 339 186 435 189
rect 339 169 345 186
rect 429 169 435 186
rect 339 166 435 169
rect -463 144 -440 150
rect -463 -144 -460 144
rect -443 -144 -440 144
rect -463 -150 -440 -144
rect -334 144 -311 150
rect -334 -144 -331 144
rect -314 -144 -311 144
rect -334 -150 -311 -144
rect -205 144 -182 150
rect -205 -144 -202 144
rect -185 -144 -182 144
rect -205 -150 -182 -144
rect -76 144 -53 150
rect -76 -144 -73 144
rect -56 -144 -53 144
rect -76 -150 -53 -144
rect 53 144 76 150
rect 53 -144 56 144
rect 73 -144 76 144
rect 53 -150 76 -144
rect 182 144 205 150
rect 182 -144 185 144
rect 202 -144 205 144
rect 182 -150 205 -144
rect 311 144 334 150
rect 311 -144 314 144
rect 331 -144 334 144
rect 311 -150 334 -144
rect 440 144 463 150
rect 440 -144 443 144
rect 460 -144 463 144
rect 440 -150 463 -144
rect -435 -169 -339 -166
rect -435 -186 -429 -169
rect -345 -186 -339 -169
rect -435 -189 -339 -186
rect -306 -169 -210 -166
rect -306 -186 -300 -169
rect -216 -186 -210 -169
rect -306 -189 -210 -186
rect -177 -169 -81 -166
rect -177 -186 -171 -169
rect -87 -186 -81 -169
rect -177 -189 -81 -186
rect -48 -169 48 -166
rect -48 -186 -42 -169
rect 42 -186 48 -169
rect -48 -189 48 -186
rect 81 -169 177 -166
rect 81 -186 87 -169
rect 171 -186 177 -169
rect 81 -189 177 -186
rect 210 -169 306 -166
rect 210 -186 216 -169
rect 300 -186 306 -169
rect 210 -189 306 -186
rect 339 -169 435 -166
rect 339 -186 345 -169
rect 429 -186 435 -169
rect 339 -189 435 -186
<< properties >>
string FIXED_BBOX -518 -246 518 246
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
