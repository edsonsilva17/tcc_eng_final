magic
tech sky130A
magscale 1 2
timestamp 1712876180
<< metal1 >>
rect 1550 14400 6680 15020
rect 1550 14280 6500 14400
rect 6620 14280 6680 14400
rect 1550 14260 6680 14280
rect 650 13110 6170 13870
rect 650 4950 810 13110
rect 1440 12980 6430 13030
rect 6270 7410 6430 12980
rect 6450 6090 6680 6290
rect 6450 5080 6680 5280
rect 630 4750 1060 4950
rect 6270 4230 6640 4250
rect 6270 4110 6500 4230
rect 6620 4110 6640 4230
rect 6270 4090 6640 4110
rect 630 3620 860 3820
<< via1 >>
rect 6500 14280 6620 14400
rect 6500 4110 6620 4230
<< metal2 >>
rect 6480 14400 6640 14420
rect 6480 14280 6500 14400
rect 6620 14280 6640 14400
rect 6480 4230 6640 14280
rect 6480 4110 6500 4230
rect 6620 4110 6640 4230
rect 6480 4090 6640 4110
use sky130_fd_pr__nfet_03v3_nvt_UUC83J  XM1
timestamp 1712876070
transform 1 0 3783 0 1 14066
box -2569 -1258 2569 1258
use Ota_esq  x1 celulas_ind
timestamp 1712866896
transform 1 0 1030 0 1 7060
box -170 -3790 5420 5650
<< labels >>
flabel metal1 630 3620 830 3820 0 FreeSans 256 0 0 0 ldo_ibias
port 4 nsew
flabel metal1 6480 6090 6680 6290 0 FreeSans 256 0 0 0 ldo_ref
port 3 nsew
flabel metal1 6480 5080 6680 5280 0 FreeSans 256 0 0 0 ldo_gnd
port 2 nsew
flabel metal1 650 13380 850 13580 0 FreeSans 256 0 0 0 ldo_in
port 1 nsew
flabel metal1 6480 14590 6680 14790 0 FreeSans 256 0 0 0 ldo_out
port 0 nsew
<< end >>
