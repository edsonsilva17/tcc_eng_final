magic
tech sky130A
magscale 1 2
timestamp 1712847951
<< metal3 >>
rect -2450 2372 2449 2400
rect -2450 -2372 2365 2372
rect 2429 -2372 2449 2372
rect -2450 -2400 2449 -2372
<< via3 >>
rect 2365 -2372 2429 2372
<< mimcap >>
rect -2350 2260 2250 2300
rect -2350 -2260 -2310 2260
rect 2210 -2260 2250 2260
rect -2350 -2300 2250 -2260
<< mimcapcontact >>
rect -2310 -2260 2210 2260
<< metal4 >>
rect 2349 2372 2445 2388
rect -2311 2260 2211 2261
rect -2311 -2260 -2310 2260
rect 2210 -2260 2211 2260
rect -2311 -2261 2211 -2260
rect 2349 -2372 2365 2372
rect 2429 -2372 2445 2372
rect 2349 -2388 2445 -2372
<< properties >>
string FIXED_BBOX -2450 -2400 2350 2400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 23.0 l 23.0 val 1.075k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
