** sch_path: /foss/designs/tcc_eng_final/xschem/multiplier-full-1-casamento-dbm.sch
**.subckt multiplier-full-1-casamento-dbm
V1 din GND sin (0 amp 2.45E9)
.save i(v1)
x1 do net3 GND cell
R2 GND do 190k m=1
R1 din net1 {Z} m=1
L3 net2 net1 2923n m=1
C2 net2 GND 0.0023393p m=1
L5 net3 net2 4710n m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt




.PARAM Z = 300
.PARAM amp = 0.24495


.CONTROL
foreach mydbm -10 -9 -8 -7 -6 -5 -4 -3 -2 -1 0
  echo amp is $mydbm
  reset
  alterparam amp = ((sqrt(2))*(sqrt(Z/1000))*(10**(($mydbm)/20)))
  save all
  tran 0.02n 5u
  meas tran out RMS v(do) from=4.999u to=5u
end

  wrdata mul1.csv tran1.out tran2.out tran3.out tran4.out tran5.out tran6.out tran7.out tran8.out
+ tran9.out tran10.out tran11.out

.ENDC

**** end user architecture code


.GLOBAL GND
.end

**** end user architecture code
**.ends

* expanding   symbol:  cell.sym # of pins=3
** sym_path: /foss/designs/tcc_eng_final/xschem/cell.sym
** sch_path: /foss/designs/tcc_eng_final/xschem/cell.sch
.subckt cell o i ground
*.iopin ground
*.iopin o
*.iopin i
XM10 net1 net1 ground net1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=40 nf=5 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 o o net1 o sky130_fd_pr__pfet_01v8_lvt L=0.35 W=40 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC3 o ground sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=3 m=3
XC2 net1 i sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=1 m=1
.ends

.GLOBAL GND
.end
