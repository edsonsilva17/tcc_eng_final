magic
tech sky130A
timestamp 1712947696
<< metal1 >>
rect 385 16560 500 16660
rect 600 16570 9755 16650
rect 385 11340 500 11440
rect 1655 11130 1750 11440
rect 4960 11430 5040 13120
rect 9530 11430 9610 13120
rect 14215 13020 14230 13120
rect 14305 13020 14320 13120
rect 17265 13020 17380 13120
rect 4960 11350 5070 11430
rect 9530 11350 9665 11430
rect 1655 11120 6415 11130
rect 1655 11040 6330 11120
rect 6405 11040 6415 11120
rect 1655 11030 6415 11040
rect 10905 11120 14445 11130
rect 10905 11040 10915 11120
rect 11005 11040 14360 11120
rect 14435 11040 14445 11120
rect 10905 11030 14445 11040
rect 17250 9355 17365 9455
rect 14240 7765 14320 7895
rect 17265 7765 17365 7775
rect 14240 7685 17365 7765
rect 17265 7675 17365 7685
<< via1 >>
rect 6330 11040 6405 11120
rect 10915 11040 11005 11120
rect 14360 11040 14435 11120
<< metal2 >>
rect 6320 11120 11015 11130
rect 6320 11040 6330 11120
rect 6405 11040 10915 11120
rect 11005 11040 11015 11120
rect 6320 11030 11015 11040
rect 14350 11120 17130 11130
rect 14350 11040 14360 11120
rect 14435 11040 17130 11120
rect 14350 11030 17130 11040
use cell  x1
timestamp 1712944235
transform 1 0 950 0 1 11250
box -450 -7700 4100 5410
use cell  x2
timestamp 1712944235
transform 1 0 5520 0 1 11250
box -450 -7700 4100 5410
use cell  x3
timestamp 1712944235
transform 1 0 10115 0 1 11250
box -450 -7700 4100 5410
use LDO  x4
timestamp 1712939325
transform 1 0 14230 0 1 7645
box 0 250 3035 5475
<< labels >>
flabel metal1 385 16560 485 16660 0 FreeSans 128 0 0 0 top_in
port 0 nsew
flabel metal1 385 11340 485 11440 0 FreeSans 128 0 0 0 top_gnd
port 1 nsew
flabel metal1 17265 7675 17365 7775 0 FreeSans 128 0 0 0 top_ibias
port 2 nsew
flabel metal1 17265 9355 17365 9455 0 FreeSans 128 0 0 0 top_ref
port 3 nsew
flabel metal1 17280 13020 17380 13120 0 FreeSans 128 0 0 0 top_out
port 4 nsew
<< end >>
