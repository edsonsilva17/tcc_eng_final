** sch_path: /foss/designs/tcc_eng_final/xschem/multiplier-full-8.sch
**.subckt multiplier-full-8
V1 in GND sin (0 1 2.45E9)
.save i(v1)
x1 net1 in GND cell
R1 out1 GND 190k m=1
x2 net2 in net1 cell
x3 net3 in net2 cell
x4 net4 in net3 cell
x5 net5 in net4 cell
x6 net6 in net5 cell
x7 net7 in net6 cell
x8 out1 in net7 cell
**** begin user architecture code


*.TRAN TSTEP TSTOP <TSTART <TMAX>> <UIC>

.control
save all
tran 0.01n 5u
wrdata ret8.csv out1
plot out1
.endc



** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  cell.sym # of pins=3
** sym_path: /foss/designs/tcc_eng_final/xschem/cell.sym
** sch_path: /foss/designs/tcc_eng_final/xschem/cell.sch
.subckt cell o i ground
*.iopin ground
*.iopin o
*.iopin i
XM10 net1 net1 ground net1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=40 nf=5 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 o o net1 o sky130_fd_pr__pfet_01v8_lvt L=0.35 W=40 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC3 o ground sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=3 m=3
XC2 net1 i sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=1 m=1
.ends

.GLOBAL GND
.end
