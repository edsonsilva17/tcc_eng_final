magic
tech sky130A
magscale 1 2
timestamp 1713011118
<< nwell >>
rect 100 16400 1074 18438
rect 1340 18000 2314 20038
rect 9230 11640 13042 12834
rect 10520 9390 13042 11640
rect 13300 10340 13916 12254
<< pwell >>
rect 11837 18901 14353 19457
rect 10842 12892 13046 14008
rect 13972 9392 14528 13208
<< nnmos >>
rect 12095 19129 14095 19229
<< mvnmos >>
rect 11070 13150 11270 13750
rect 11328 13150 11528 13750
rect 11586 13150 11786 13750
rect 11844 13150 12044 13750
rect 12102 13150 12302 13750
rect 12360 13150 12560 13750
rect 12618 13150 12818 13750
rect 14200 11550 14300 12950
rect 14200 9650 14300 11050
<< mvpmos >>
rect 9488 11937 9688 12537
rect 9746 11937 9946 12537
rect 10004 11937 10204 12537
rect 10262 11937 10462 12537
rect 10520 11937 10720 12537
rect 10778 11937 10978 12537
rect 11036 11937 11236 12537
rect 11294 11937 11494 12537
rect 11552 11937 11752 12537
rect 11810 11937 12010 12537
rect 12068 11937 12268 12537
rect 12326 11937 12526 12537
rect 12584 11937 12784 12537
rect 10778 10817 10978 11417
rect 11036 10817 11236 11417
rect 11294 10817 11494 11417
rect 11552 10817 11752 11417
rect 11810 10817 12010 11417
rect 12068 10817 12268 11417
rect 12326 10817 12526 11417
rect 12584 10817 12784 11417
rect 13558 11557 13658 11957
rect 10778 9687 10978 10287
rect 11036 9687 11236 10287
rect 11294 9687 11494 10287
rect 11552 9687 11752 10287
rect 11810 9687 12010 10287
rect 12068 9687 12268 10287
rect 12326 9687 12526 10287
rect 12584 9687 12784 10287
rect 13558 10637 13658 11037
<< pmoslvt >>
rect 296 16619 366 18219
rect 424 16619 494 18219
rect 552 16619 622 18219
rect 680 16619 750 18219
rect 808 16619 878 18219
rect 1536 18219 1606 19819
rect 1664 18219 1734 19819
rect 1792 18219 1862 19819
rect 1920 18219 1990 19819
rect 2048 18219 2118 19819
<< pdiff >>
rect 238 18207 296 18219
rect 238 16631 250 18207
rect 284 16631 296 18207
rect 238 16619 296 16631
rect 366 18207 424 18219
rect 366 16631 378 18207
rect 412 16631 424 18207
rect 366 16619 424 16631
rect 494 18207 552 18219
rect 494 16631 506 18207
rect 540 16631 552 18207
rect 494 16619 552 16631
rect 622 18207 680 18219
rect 622 16631 634 18207
rect 668 16631 680 18207
rect 622 16619 680 16631
rect 750 18207 808 18219
rect 750 16631 762 18207
rect 796 16631 808 18207
rect 750 16619 808 16631
rect 878 18207 936 18219
rect 878 16631 890 18207
rect 924 16631 936 18207
rect 878 16619 936 16631
rect 1478 19807 1536 19819
rect 1478 18231 1490 19807
rect 1524 18231 1536 19807
rect 1478 18219 1536 18231
rect 1606 19807 1664 19819
rect 1606 18231 1618 19807
rect 1652 18231 1664 19807
rect 1606 18219 1664 18231
rect 1734 19807 1792 19819
rect 1734 18231 1746 19807
rect 1780 18231 1792 19807
rect 1734 18219 1792 18231
rect 1862 19807 1920 19819
rect 1862 18231 1874 19807
rect 1908 18231 1920 19807
rect 1862 18219 1920 18231
rect 1990 19807 2048 19819
rect 1990 18231 2002 19807
rect 2036 18231 2048 19807
rect 1990 18219 2048 18231
rect 2118 19807 2176 19819
rect 2118 18231 2130 19807
rect 2164 18231 2176 19807
rect 2118 18219 2176 18231
<< mvndiff >>
rect 12095 19275 14095 19287
rect 12095 19241 12107 19275
rect 14083 19241 14095 19275
rect 12095 19229 14095 19241
rect 12095 19117 14095 19129
rect 12095 19083 12107 19117
rect 14083 19083 14095 19117
rect 12095 19071 14095 19083
rect 11012 13738 11070 13750
rect 11012 13162 11024 13738
rect 11058 13162 11070 13738
rect 11012 13150 11070 13162
rect 11270 13738 11328 13750
rect 11270 13162 11282 13738
rect 11316 13162 11328 13738
rect 11270 13150 11328 13162
rect 11528 13738 11586 13750
rect 11528 13162 11540 13738
rect 11574 13162 11586 13738
rect 11528 13150 11586 13162
rect 11786 13738 11844 13750
rect 11786 13162 11798 13738
rect 11832 13162 11844 13738
rect 11786 13150 11844 13162
rect 12044 13738 12102 13750
rect 12044 13162 12056 13738
rect 12090 13162 12102 13738
rect 12044 13150 12102 13162
rect 12302 13738 12360 13750
rect 12302 13162 12314 13738
rect 12348 13162 12360 13738
rect 12302 13150 12360 13162
rect 12560 13738 12618 13750
rect 12560 13162 12572 13738
rect 12606 13162 12618 13738
rect 12560 13150 12618 13162
rect 12818 13738 12876 13750
rect 12818 13162 12830 13738
rect 12864 13162 12876 13738
rect 12818 13150 12876 13162
rect 14142 12938 14200 12950
rect 14142 11562 14154 12938
rect 14188 11562 14200 12938
rect 14142 11550 14200 11562
rect 14300 12938 14358 12950
rect 14300 11562 14312 12938
rect 14346 11562 14358 12938
rect 14300 11550 14358 11562
rect 14142 11038 14200 11050
rect 14142 9662 14154 11038
rect 14188 9662 14200 11038
rect 14142 9650 14200 9662
rect 14300 11038 14358 11050
rect 14300 9662 14312 11038
rect 14346 9662 14358 11038
rect 14300 9650 14358 9662
<< mvpdiff >>
rect 9430 12525 9488 12537
rect 9430 11949 9442 12525
rect 9476 11949 9488 12525
rect 9430 11937 9488 11949
rect 9688 12525 9746 12537
rect 9688 11949 9700 12525
rect 9734 11949 9746 12525
rect 9688 11937 9746 11949
rect 9946 12525 10004 12537
rect 9946 11949 9958 12525
rect 9992 11949 10004 12525
rect 9946 11937 10004 11949
rect 10204 12525 10262 12537
rect 10204 11949 10216 12525
rect 10250 11949 10262 12525
rect 10204 11937 10262 11949
rect 10462 12525 10520 12537
rect 10462 11949 10474 12525
rect 10508 11949 10520 12525
rect 10462 11937 10520 11949
rect 10720 12525 10778 12537
rect 10720 11949 10732 12525
rect 10766 11949 10778 12525
rect 10720 11937 10778 11949
rect 10978 12525 11036 12537
rect 10978 11949 10990 12525
rect 11024 11949 11036 12525
rect 10978 11937 11036 11949
rect 11236 12525 11294 12537
rect 11236 11949 11248 12525
rect 11282 11949 11294 12525
rect 11236 11937 11294 11949
rect 11494 12525 11552 12537
rect 11494 11949 11506 12525
rect 11540 11949 11552 12525
rect 11494 11937 11552 11949
rect 11752 12525 11810 12537
rect 11752 11949 11764 12525
rect 11798 11949 11810 12525
rect 11752 11937 11810 11949
rect 12010 12525 12068 12537
rect 12010 11949 12022 12525
rect 12056 11949 12068 12525
rect 12010 11937 12068 11949
rect 12268 12525 12326 12537
rect 12268 11949 12280 12525
rect 12314 11949 12326 12525
rect 12268 11937 12326 11949
rect 12526 12525 12584 12537
rect 12526 11949 12538 12525
rect 12572 11949 12584 12525
rect 12526 11937 12584 11949
rect 12784 12525 12842 12537
rect 12784 11949 12796 12525
rect 12830 11949 12842 12525
rect 12784 11937 12842 11949
rect 10720 11405 10778 11417
rect 10720 10829 10732 11405
rect 10766 10829 10778 11405
rect 10720 10817 10778 10829
rect 10978 11405 11036 11417
rect 10978 10829 10990 11405
rect 11024 10829 11036 11405
rect 10978 10817 11036 10829
rect 11236 11405 11294 11417
rect 11236 10829 11248 11405
rect 11282 10829 11294 11405
rect 11236 10817 11294 10829
rect 11494 11405 11552 11417
rect 11494 10829 11506 11405
rect 11540 10829 11552 11405
rect 11494 10817 11552 10829
rect 11752 11405 11810 11417
rect 11752 10829 11764 11405
rect 11798 10829 11810 11405
rect 11752 10817 11810 10829
rect 12010 11405 12068 11417
rect 12010 10829 12022 11405
rect 12056 10829 12068 11405
rect 12010 10817 12068 10829
rect 12268 11405 12326 11417
rect 12268 10829 12280 11405
rect 12314 10829 12326 11405
rect 12268 10817 12326 10829
rect 12526 11405 12584 11417
rect 12526 10829 12538 11405
rect 12572 10829 12584 11405
rect 12526 10817 12584 10829
rect 12784 11405 12842 11417
rect 12784 10829 12796 11405
rect 12830 10829 12842 11405
rect 12784 10817 12842 10829
rect 13500 11945 13558 11957
rect 13500 11569 13512 11945
rect 13546 11569 13558 11945
rect 13500 11557 13558 11569
rect 13658 11945 13716 11957
rect 13658 11569 13670 11945
rect 13704 11569 13716 11945
rect 13658 11557 13716 11569
rect 10720 10275 10778 10287
rect 10720 9699 10732 10275
rect 10766 9699 10778 10275
rect 10720 9687 10778 9699
rect 10978 10275 11036 10287
rect 10978 9699 10990 10275
rect 11024 9699 11036 10275
rect 10978 9687 11036 9699
rect 11236 10275 11294 10287
rect 11236 9699 11248 10275
rect 11282 9699 11294 10275
rect 11236 9687 11294 9699
rect 11494 10275 11552 10287
rect 11494 9699 11506 10275
rect 11540 9699 11552 10275
rect 11494 9687 11552 9699
rect 11752 10275 11810 10287
rect 11752 9699 11764 10275
rect 11798 9699 11810 10275
rect 11752 9687 11810 9699
rect 12010 10275 12068 10287
rect 12010 9699 12022 10275
rect 12056 9699 12068 10275
rect 12010 9687 12068 9699
rect 12268 10275 12326 10287
rect 12268 9699 12280 10275
rect 12314 9699 12326 10275
rect 12268 9687 12326 9699
rect 12526 10275 12584 10287
rect 12526 9699 12538 10275
rect 12572 9699 12584 10275
rect 12526 9687 12584 9699
rect 12784 10275 12842 10287
rect 12784 9699 12796 10275
rect 12830 9699 12842 10275
rect 12784 9687 12842 9699
rect 13500 11025 13558 11037
rect 13500 10649 13512 11025
rect 13546 10649 13558 11025
rect 13500 10637 13558 10649
rect 13658 11025 13716 11037
rect 13658 10649 13670 11025
rect 13704 10649 13716 11025
rect 13658 10637 13716 10649
<< pdiffc >>
rect 250 16631 284 18207
rect 378 16631 412 18207
rect 506 16631 540 18207
rect 634 16631 668 18207
rect 762 16631 796 18207
rect 890 16631 924 18207
rect 1490 18231 1524 19807
rect 1618 18231 1652 19807
rect 1746 18231 1780 19807
rect 1874 18231 1908 19807
rect 2002 18231 2036 19807
rect 2130 18231 2164 19807
<< mvndiffc >>
rect 12107 19241 14083 19275
rect 12107 19083 14083 19117
rect 11024 13162 11058 13738
rect 11282 13162 11316 13738
rect 11540 13162 11574 13738
rect 11798 13162 11832 13738
rect 12056 13162 12090 13738
rect 12314 13162 12348 13738
rect 12572 13162 12606 13738
rect 12830 13162 12864 13738
rect 14154 11562 14188 12938
rect 14312 11562 14346 12938
rect 14154 9662 14188 11038
rect 14312 9662 14346 11038
<< mvpdiffc >>
rect 9442 11949 9476 12525
rect 9700 11949 9734 12525
rect 9958 11949 9992 12525
rect 10216 11949 10250 12525
rect 10474 11949 10508 12525
rect 10732 11949 10766 12525
rect 10990 11949 11024 12525
rect 11248 11949 11282 12525
rect 11506 11949 11540 12525
rect 11764 11949 11798 12525
rect 12022 11949 12056 12525
rect 12280 11949 12314 12525
rect 12538 11949 12572 12525
rect 12796 11949 12830 12525
rect 10732 10829 10766 11405
rect 10990 10829 11024 11405
rect 11248 10829 11282 11405
rect 11506 10829 11540 11405
rect 11764 10829 11798 11405
rect 12022 10829 12056 11405
rect 12280 10829 12314 11405
rect 12538 10829 12572 11405
rect 12796 10829 12830 11405
rect 13512 11569 13546 11945
rect 13670 11569 13704 11945
rect 10732 9699 10766 10275
rect 10990 9699 11024 10275
rect 11248 9699 11282 10275
rect 11506 9699 11540 10275
rect 11764 9699 11798 10275
rect 12022 9699 12056 10275
rect 12280 9699 12314 10275
rect 12538 9699 12572 10275
rect 12796 9699 12830 10275
rect 13512 10649 13546 11025
rect 13670 10649 13704 11025
<< nsubdiff >>
rect 1376 19968 1472 20002
rect 2182 19968 2278 20002
rect 1376 19906 1410 19968
rect 136 18368 232 18402
rect 942 18368 1038 18402
rect 136 18306 170 18368
rect 1004 18306 1038 18368
rect 136 16470 170 16532
rect 2244 19906 2278 19968
rect 1376 18070 1410 18132
rect 2244 18070 2278 18132
rect 1376 18036 1472 18070
rect 2182 18036 2278 18070
rect 1004 16470 1038 16532
rect 136 16436 232 16470
rect 942 16436 1038 16470
<< mvpsubdiff >>
rect 11873 19409 14317 19421
rect 11873 19375 11981 19409
rect 14209 19375 14317 19409
rect 11873 19363 14317 19375
rect 11873 19313 11931 19363
rect 11873 19045 11885 19313
rect 11919 19045 11931 19313
rect 14259 19313 14317 19363
rect 11873 18995 11931 19045
rect 14259 19045 14271 19313
rect 14305 19045 14317 19313
rect 14259 18995 14317 19045
rect 11873 18983 14317 18995
rect 11873 18949 11981 18983
rect 14209 18949 14317 18983
rect 11873 18937 14317 18949
rect 10878 13960 13010 13972
rect 10878 13926 10986 13960
rect 12902 13926 13010 13960
rect 10878 13914 13010 13926
rect 10878 13864 10936 13914
rect 10878 13036 10890 13864
rect 10924 13036 10936 13864
rect 12952 13864 13010 13914
rect 10878 12986 10936 13036
rect 12952 13036 12964 13864
rect 12998 13036 13010 13864
rect 12952 12986 13010 13036
rect 10878 12974 13010 12986
rect 10878 12940 10986 12974
rect 12902 12940 13010 12974
rect 10878 12928 13010 12940
rect 14008 13160 14492 13172
rect 14008 13126 14116 13160
rect 14384 13126 14492 13160
rect 14008 13114 14492 13126
rect 14008 13064 14066 13114
rect 14008 11436 14020 13064
rect 14054 11436 14066 13064
rect 14434 13064 14492 13114
rect 14008 11386 14066 11436
rect 14434 11436 14446 13064
rect 14480 11436 14492 13064
rect 14434 11386 14492 11436
rect 14008 11374 14492 11386
rect 14008 11340 14116 11374
rect 14384 11340 14492 11374
rect 14008 11328 14492 11340
rect 14008 11260 14492 11272
rect 14008 11226 14116 11260
rect 14384 11226 14492 11260
rect 14008 11214 14492 11226
rect 14008 11164 14066 11214
rect 14008 9536 14020 11164
rect 14054 9536 14066 11164
rect 14434 11164 14492 11214
rect 14008 9486 14066 9536
rect 14434 9536 14446 11164
rect 14480 9536 14492 11164
rect 14434 9486 14492 9536
rect 14008 9474 14492 9486
rect 14008 9440 14116 9474
rect 14384 9440 14492 9474
rect 14008 9428 14492 9440
<< mvnsubdiff >>
rect 9296 12756 12976 12768
rect 9296 12722 9404 12756
rect 12868 12722 12976 12756
rect 9296 12710 12976 12722
rect 9296 12660 9354 12710
rect 9296 11814 9308 12660
rect 9342 11814 9354 12660
rect 12918 12660 12976 12710
rect 9296 11764 9354 11814
rect 12918 11814 12930 12660
rect 12964 11814 12976 12660
rect 12918 11764 12976 11814
rect 9296 11752 12976 11764
rect 9296 11718 9404 11752
rect 12868 11718 12976 11752
rect 9296 11706 12976 11718
rect 13366 12176 13850 12188
rect 13366 12142 13474 12176
rect 13742 12142 13850 12176
rect 13366 12130 13850 12142
rect 13366 12080 13424 12130
rect 10586 11636 12976 11648
rect 10586 11602 10694 11636
rect 12868 11602 12976 11636
rect 10586 11590 12976 11602
rect 10586 11540 10644 11590
rect 10586 10694 10598 11540
rect 10632 10694 10644 11540
rect 12918 11540 12976 11590
rect 10586 10644 10644 10694
rect 12918 10694 12930 11540
rect 12964 10694 12976 11540
rect 13366 11434 13378 12080
rect 13412 11434 13424 12080
rect 13792 12080 13850 12130
rect 13366 11384 13424 11434
rect 13792 11434 13804 12080
rect 13838 11434 13850 12080
rect 13792 11384 13850 11434
rect 13366 11372 13850 11384
rect 13366 11338 13474 11372
rect 13742 11338 13850 11372
rect 13366 11326 13850 11338
rect 12918 10644 12976 10694
rect 10586 10632 12976 10644
rect 10586 10598 10694 10632
rect 12868 10598 12976 10632
rect 10586 10586 12976 10598
rect 13366 11256 13850 11268
rect 13366 11222 13474 11256
rect 13742 11222 13850 11256
rect 13366 11210 13850 11222
rect 13366 11160 13424 11210
rect 10586 10506 12976 10518
rect 10586 10472 10694 10506
rect 12868 10472 12976 10506
rect 10586 10460 12976 10472
rect 10586 10410 10644 10460
rect 10586 9564 10598 10410
rect 10632 9564 10644 10410
rect 12918 10410 12976 10460
rect 10586 9514 10644 9564
rect 12918 9564 12930 10410
rect 12964 9564 12976 10410
rect 13366 10514 13378 11160
rect 13412 10514 13424 11160
rect 13792 11160 13850 11210
rect 13366 10464 13424 10514
rect 13792 10514 13804 11160
rect 13838 10514 13850 11160
rect 13792 10464 13850 10514
rect 13366 10452 13850 10464
rect 13366 10418 13474 10452
rect 13742 10418 13850 10452
rect 13366 10406 13850 10418
rect 12918 9514 12976 9564
rect 10586 9502 12976 9514
rect 10586 9468 10694 9502
rect 12868 9468 12976 9502
rect 10586 9456 12976 9468
<< nsubdiffcont >>
rect 1472 19968 2182 20002
rect 232 18368 942 18402
rect 136 16532 170 18306
rect 1004 16532 1038 18306
rect 1376 18132 1410 19906
rect 2244 18132 2278 19906
rect 1472 18036 2182 18070
rect 232 16436 942 16470
<< mvpsubdiffcont >>
rect 11981 19375 14209 19409
rect 11885 19045 11919 19313
rect 14271 19045 14305 19313
rect 11981 18949 14209 18983
rect 10986 13926 12902 13960
rect 10890 13036 10924 13864
rect 12964 13036 12998 13864
rect 10986 12940 12902 12974
rect 14116 13126 14384 13160
rect 14020 11436 14054 13064
rect 14446 11436 14480 13064
rect 14116 11340 14384 11374
rect 14116 11226 14384 11260
rect 14020 9536 14054 11164
rect 14446 9536 14480 11164
rect 14116 9440 14384 9474
<< mvnsubdiffcont >>
rect 9404 12722 12868 12756
rect 9308 11814 9342 12660
rect 12930 11814 12964 12660
rect 9404 11718 12868 11752
rect 13474 12142 13742 12176
rect 10694 11602 12868 11636
rect 10598 10694 10632 11540
rect 12930 10694 12964 11540
rect 13378 11434 13412 12080
rect 13804 11434 13838 12080
rect 13474 11338 13742 11372
rect 10694 10598 12868 10632
rect 13474 11222 13742 11256
rect 10694 10472 12868 10506
rect 10598 9564 10632 10410
rect 12930 9564 12964 10410
rect 13378 10514 13412 11160
rect 13804 10514 13838 11160
rect 13474 10418 13742 10452
rect 10694 9468 12868 9502
<< poly >>
rect 296 18300 366 18316
rect 296 18266 312 18300
rect 350 18266 366 18300
rect 296 18219 366 18266
rect 424 18300 494 18316
rect 424 18266 440 18300
rect 478 18266 494 18300
rect 424 18219 494 18266
rect 552 18300 622 18316
rect 552 18266 568 18300
rect 606 18266 622 18300
rect 552 18219 622 18266
rect 680 18300 750 18316
rect 680 18266 696 18300
rect 734 18266 750 18300
rect 680 18219 750 18266
rect 808 18300 878 18316
rect 808 18266 824 18300
rect 862 18266 878 18300
rect 808 18219 878 18266
rect 296 16572 366 16619
rect 296 16538 312 16572
rect 350 16538 366 16572
rect 296 16522 366 16538
rect 424 16572 494 16619
rect 424 16538 440 16572
rect 478 16538 494 16572
rect 424 16522 494 16538
rect 552 16572 622 16619
rect 552 16538 568 16572
rect 606 16538 622 16572
rect 552 16522 622 16538
rect 680 16572 750 16619
rect 680 16538 696 16572
rect 734 16538 750 16572
rect 680 16522 750 16538
rect 808 16572 878 16619
rect 808 16538 824 16572
rect 862 16538 878 16572
rect 808 16522 878 16538
rect 1536 19900 1606 19916
rect 1536 19866 1552 19900
rect 1590 19866 1606 19900
rect 1536 19819 1606 19866
rect 1664 19900 1734 19916
rect 1664 19866 1680 19900
rect 1718 19866 1734 19900
rect 1664 19819 1734 19866
rect 1792 19900 1862 19916
rect 1792 19866 1808 19900
rect 1846 19866 1862 19900
rect 1792 19819 1862 19866
rect 1920 19900 1990 19916
rect 1920 19866 1936 19900
rect 1974 19866 1990 19900
rect 1920 19819 1990 19866
rect 2048 19900 2118 19916
rect 2048 19866 2064 19900
rect 2102 19866 2118 19900
rect 2048 19819 2118 19866
rect 1536 18172 1606 18219
rect 1536 18138 1552 18172
rect 1590 18138 1606 18172
rect 1536 18122 1606 18138
rect 1664 18172 1734 18219
rect 1664 18138 1680 18172
rect 1718 18138 1734 18172
rect 1664 18122 1734 18138
rect 1792 18172 1862 18219
rect 1792 18138 1808 18172
rect 1846 18138 1862 18172
rect 1792 18122 1862 18138
rect 1920 18172 1990 18219
rect 1920 18138 1936 18172
rect 1974 18138 1990 18172
rect 1920 18122 1990 18138
rect 2048 18172 2118 18219
rect 2048 18138 2064 18172
rect 2102 18138 2118 18172
rect 2048 18122 2118 18138
rect 12007 19213 12095 19229
rect 12007 19145 12023 19213
rect 12057 19145 12095 19213
rect 12007 19129 12095 19145
rect 14095 19213 14183 19229
rect 14095 19145 14133 19213
rect 14167 19145 14183 19213
rect 14095 19129 14183 19145
rect 11070 13822 11270 13838
rect 11070 13788 11086 13822
rect 11254 13788 11270 13822
rect 11070 13750 11270 13788
rect 11328 13822 11528 13838
rect 11328 13788 11344 13822
rect 11512 13788 11528 13822
rect 11328 13750 11528 13788
rect 11586 13822 11786 13838
rect 11586 13788 11602 13822
rect 11770 13788 11786 13822
rect 11586 13750 11786 13788
rect 11844 13822 12044 13838
rect 11844 13788 11860 13822
rect 12028 13788 12044 13822
rect 11844 13750 12044 13788
rect 12102 13822 12302 13838
rect 12102 13788 12118 13822
rect 12286 13788 12302 13822
rect 12102 13750 12302 13788
rect 12360 13822 12560 13838
rect 12360 13788 12376 13822
rect 12544 13788 12560 13822
rect 12360 13750 12560 13788
rect 12618 13822 12818 13838
rect 12618 13788 12634 13822
rect 12802 13788 12818 13822
rect 12618 13750 12818 13788
rect 11070 13112 11270 13150
rect 11070 13078 11086 13112
rect 11254 13078 11270 13112
rect 11070 13062 11270 13078
rect 11328 13112 11528 13150
rect 11328 13078 11344 13112
rect 11512 13078 11528 13112
rect 11328 13062 11528 13078
rect 11586 13112 11786 13150
rect 11586 13078 11602 13112
rect 11770 13078 11786 13112
rect 11586 13062 11786 13078
rect 11844 13112 12044 13150
rect 11844 13078 11860 13112
rect 12028 13078 12044 13112
rect 11844 13062 12044 13078
rect 12102 13112 12302 13150
rect 12102 13078 12118 13112
rect 12286 13078 12302 13112
rect 12102 13062 12302 13078
rect 12360 13112 12560 13150
rect 12360 13078 12376 13112
rect 12544 13078 12560 13112
rect 12360 13062 12560 13078
rect 12618 13112 12818 13150
rect 12618 13078 12634 13112
rect 12802 13078 12818 13112
rect 12618 13062 12818 13078
rect 9488 12618 9688 12634
rect 9488 12584 9504 12618
rect 9672 12584 9688 12618
rect 9488 12537 9688 12584
rect 9746 12618 9946 12634
rect 9746 12584 9762 12618
rect 9930 12584 9946 12618
rect 9746 12537 9946 12584
rect 10004 12618 10204 12634
rect 10004 12584 10020 12618
rect 10188 12584 10204 12618
rect 10004 12537 10204 12584
rect 10262 12618 10462 12634
rect 10262 12584 10278 12618
rect 10446 12584 10462 12618
rect 10262 12537 10462 12584
rect 10520 12618 10720 12634
rect 10520 12584 10536 12618
rect 10704 12584 10720 12618
rect 10520 12537 10720 12584
rect 10778 12618 10978 12634
rect 10778 12584 10794 12618
rect 10962 12584 10978 12618
rect 10778 12537 10978 12584
rect 11036 12618 11236 12634
rect 11036 12584 11052 12618
rect 11220 12584 11236 12618
rect 11036 12537 11236 12584
rect 11294 12618 11494 12634
rect 11294 12584 11310 12618
rect 11478 12584 11494 12618
rect 11294 12537 11494 12584
rect 11552 12618 11752 12634
rect 11552 12584 11568 12618
rect 11736 12584 11752 12618
rect 11552 12537 11752 12584
rect 11810 12618 12010 12634
rect 11810 12584 11826 12618
rect 11994 12584 12010 12618
rect 11810 12537 12010 12584
rect 12068 12618 12268 12634
rect 12068 12584 12084 12618
rect 12252 12584 12268 12618
rect 12068 12537 12268 12584
rect 12326 12618 12526 12634
rect 12326 12584 12342 12618
rect 12510 12584 12526 12618
rect 12326 12537 12526 12584
rect 12584 12618 12784 12634
rect 12584 12584 12600 12618
rect 12768 12584 12784 12618
rect 12584 12537 12784 12584
rect 9488 11890 9688 11937
rect 9488 11856 9504 11890
rect 9672 11856 9688 11890
rect 9488 11840 9688 11856
rect 9746 11890 9946 11937
rect 9746 11856 9762 11890
rect 9930 11856 9946 11890
rect 9746 11840 9946 11856
rect 10004 11890 10204 11937
rect 10004 11856 10020 11890
rect 10188 11856 10204 11890
rect 10004 11840 10204 11856
rect 10262 11890 10462 11937
rect 10262 11856 10278 11890
rect 10446 11856 10462 11890
rect 10262 11840 10462 11856
rect 10520 11890 10720 11937
rect 10520 11856 10536 11890
rect 10704 11856 10720 11890
rect 10520 11840 10720 11856
rect 10778 11890 10978 11937
rect 10778 11856 10794 11890
rect 10962 11856 10978 11890
rect 10778 11840 10978 11856
rect 11036 11890 11236 11937
rect 11036 11856 11052 11890
rect 11220 11856 11236 11890
rect 11036 11840 11236 11856
rect 11294 11890 11494 11937
rect 11294 11856 11310 11890
rect 11478 11856 11494 11890
rect 11294 11840 11494 11856
rect 11552 11890 11752 11937
rect 11552 11856 11568 11890
rect 11736 11856 11752 11890
rect 11552 11840 11752 11856
rect 11810 11890 12010 11937
rect 11810 11856 11826 11890
rect 11994 11856 12010 11890
rect 11810 11840 12010 11856
rect 12068 11890 12268 11937
rect 12068 11856 12084 11890
rect 12252 11856 12268 11890
rect 12068 11840 12268 11856
rect 12326 11890 12526 11937
rect 12326 11856 12342 11890
rect 12510 11856 12526 11890
rect 12326 11840 12526 11856
rect 12584 11890 12784 11937
rect 12584 11856 12600 11890
rect 12768 11856 12784 11890
rect 12584 11840 12784 11856
rect 10778 11498 10978 11514
rect 10778 11464 10794 11498
rect 10962 11464 10978 11498
rect 10778 11417 10978 11464
rect 11036 11498 11236 11514
rect 11036 11464 11052 11498
rect 11220 11464 11236 11498
rect 11036 11417 11236 11464
rect 11294 11498 11494 11514
rect 11294 11464 11310 11498
rect 11478 11464 11494 11498
rect 11294 11417 11494 11464
rect 11552 11498 11752 11514
rect 11552 11464 11568 11498
rect 11736 11464 11752 11498
rect 11552 11417 11752 11464
rect 11810 11498 12010 11514
rect 11810 11464 11826 11498
rect 11994 11464 12010 11498
rect 11810 11417 12010 11464
rect 12068 11498 12268 11514
rect 12068 11464 12084 11498
rect 12252 11464 12268 11498
rect 12068 11417 12268 11464
rect 12326 11498 12526 11514
rect 12326 11464 12342 11498
rect 12510 11464 12526 11498
rect 12326 11417 12526 11464
rect 12584 11498 12784 11514
rect 12584 11464 12600 11498
rect 12768 11464 12784 11498
rect 12584 11417 12784 11464
rect 10778 10770 10978 10817
rect 10778 10736 10794 10770
rect 10962 10736 10978 10770
rect 10778 10720 10978 10736
rect 11036 10770 11236 10817
rect 11036 10736 11052 10770
rect 11220 10736 11236 10770
rect 11036 10720 11236 10736
rect 11294 10770 11494 10817
rect 11294 10736 11310 10770
rect 11478 10736 11494 10770
rect 11294 10720 11494 10736
rect 11552 10770 11752 10817
rect 11552 10736 11568 10770
rect 11736 10736 11752 10770
rect 11552 10720 11752 10736
rect 11810 10770 12010 10817
rect 11810 10736 11826 10770
rect 11994 10736 12010 10770
rect 11810 10720 12010 10736
rect 12068 10770 12268 10817
rect 12068 10736 12084 10770
rect 12252 10736 12268 10770
rect 12068 10720 12268 10736
rect 12326 10770 12526 10817
rect 12326 10736 12342 10770
rect 12510 10736 12526 10770
rect 12326 10720 12526 10736
rect 12584 10770 12784 10817
rect 12584 10736 12600 10770
rect 12768 10736 12784 10770
rect 12584 10720 12784 10736
rect 13558 12038 13658 12054
rect 13558 12004 13574 12038
rect 13642 12004 13658 12038
rect 13558 11957 13658 12004
rect 13558 11510 13658 11557
rect 13558 11476 13574 11510
rect 13642 11476 13658 11510
rect 13558 11460 13658 11476
rect 14200 13022 14300 13038
rect 14200 12988 14216 13022
rect 14284 12988 14300 13022
rect 14200 12950 14300 12988
rect 14200 11512 14300 11550
rect 14200 11478 14216 11512
rect 14284 11478 14300 11512
rect 14200 11462 14300 11478
rect 10778 10368 10978 10384
rect 10778 10334 10794 10368
rect 10962 10334 10978 10368
rect 10778 10287 10978 10334
rect 11036 10368 11236 10384
rect 11036 10334 11052 10368
rect 11220 10334 11236 10368
rect 11036 10287 11236 10334
rect 11294 10368 11494 10384
rect 11294 10334 11310 10368
rect 11478 10334 11494 10368
rect 11294 10287 11494 10334
rect 11552 10368 11752 10384
rect 11552 10334 11568 10368
rect 11736 10334 11752 10368
rect 11552 10287 11752 10334
rect 11810 10368 12010 10384
rect 11810 10334 11826 10368
rect 11994 10334 12010 10368
rect 11810 10287 12010 10334
rect 12068 10368 12268 10384
rect 12068 10334 12084 10368
rect 12252 10334 12268 10368
rect 12068 10287 12268 10334
rect 12326 10368 12526 10384
rect 12326 10334 12342 10368
rect 12510 10334 12526 10368
rect 12326 10287 12526 10334
rect 12584 10368 12784 10384
rect 12584 10334 12600 10368
rect 12768 10334 12784 10368
rect 12584 10287 12784 10334
rect 10778 9640 10978 9687
rect 10778 9606 10794 9640
rect 10962 9606 10978 9640
rect 10778 9590 10978 9606
rect 11036 9640 11236 9687
rect 11036 9606 11052 9640
rect 11220 9606 11236 9640
rect 11036 9590 11236 9606
rect 11294 9640 11494 9687
rect 11294 9606 11310 9640
rect 11478 9606 11494 9640
rect 11294 9590 11494 9606
rect 11552 9640 11752 9687
rect 11552 9606 11568 9640
rect 11736 9606 11752 9640
rect 11552 9590 11752 9606
rect 11810 9640 12010 9687
rect 11810 9606 11826 9640
rect 11994 9606 12010 9640
rect 11810 9590 12010 9606
rect 12068 9640 12268 9687
rect 12068 9606 12084 9640
rect 12252 9606 12268 9640
rect 12068 9590 12268 9606
rect 12326 9640 12526 9687
rect 12326 9606 12342 9640
rect 12510 9606 12526 9640
rect 12326 9590 12526 9606
rect 12584 9640 12784 9687
rect 12584 9606 12600 9640
rect 12768 9606 12784 9640
rect 12584 9590 12784 9606
rect 13558 11118 13658 11134
rect 13558 11084 13574 11118
rect 13642 11084 13658 11118
rect 13558 11037 13658 11084
rect 13558 10590 13658 10637
rect 13558 10556 13574 10590
rect 13642 10556 13658 10590
rect 13558 10540 13658 10556
rect 14200 11122 14300 11138
rect 14200 11088 14216 11122
rect 14284 11088 14300 11122
rect 14200 11050 14300 11088
rect 14200 9612 14300 9650
rect 14200 9578 14216 9612
rect 14284 9578 14300 9612
rect 14200 9562 14300 9578
<< polycont >>
rect 312 18266 350 18300
rect 440 18266 478 18300
rect 568 18266 606 18300
rect 696 18266 734 18300
rect 824 18266 862 18300
rect 312 16538 350 16572
rect 440 16538 478 16572
rect 568 16538 606 16572
rect 696 16538 734 16572
rect 824 16538 862 16572
rect 1552 19866 1590 19900
rect 1680 19866 1718 19900
rect 1808 19866 1846 19900
rect 1936 19866 1974 19900
rect 2064 19866 2102 19900
rect 1552 18138 1590 18172
rect 1680 18138 1718 18172
rect 1808 18138 1846 18172
rect 1936 18138 1974 18172
rect 2064 18138 2102 18172
rect 12023 19145 12057 19213
rect 14133 19145 14167 19213
rect 11086 13788 11254 13822
rect 11344 13788 11512 13822
rect 11602 13788 11770 13822
rect 11860 13788 12028 13822
rect 12118 13788 12286 13822
rect 12376 13788 12544 13822
rect 12634 13788 12802 13822
rect 11086 13078 11254 13112
rect 11344 13078 11512 13112
rect 11602 13078 11770 13112
rect 11860 13078 12028 13112
rect 12118 13078 12286 13112
rect 12376 13078 12544 13112
rect 12634 13078 12802 13112
rect 9504 12584 9672 12618
rect 9762 12584 9930 12618
rect 10020 12584 10188 12618
rect 10278 12584 10446 12618
rect 10536 12584 10704 12618
rect 10794 12584 10962 12618
rect 11052 12584 11220 12618
rect 11310 12584 11478 12618
rect 11568 12584 11736 12618
rect 11826 12584 11994 12618
rect 12084 12584 12252 12618
rect 12342 12584 12510 12618
rect 12600 12584 12768 12618
rect 9504 11856 9672 11890
rect 9762 11856 9930 11890
rect 10020 11856 10188 11890
rect 10278 11856 10446 11890
rect 10536 11856 10704 11890
rect 10794 11856 10962 11890
rect 11052 11856 11220 11890
rect 11310 11856 11478 11890
rect 11568 11856 11736 11890
rect 11826 11856 11994 11890
rect 12084 11856 12252 11890
rect 12342 11856 12510 11890
rect 12600 11856 12768 11890
rect 10794 11464 10962 11498
rect 11052 11464 11220 11498
rect 11310 11464 11478 11498
rect 11568 11464 11736 11498
rect 11826 11464 11994 11498
rect 12084 11464 12252 11498
rect 12342 11464 12510 11498
rect 12600 11464 12768 11498
rect 10794 10736 10962 10770
rect 11052 10736 11220 10770
rect 11310 10736 11478 10770
rect 11568 10736 11736 10770
rect 11826 10736 11994 10770
rect 12084 10736 12252 10770
rect 12342 10736 12510 10770
rect 12600 10736 12768 10770
rect 13574 12004 13642 12038
rect 13574 11476 13642 11510
rect 14216 12988 14284 13022
rect 14216 11478 14284 11512
rect 10794 10334 10962 10368
rect 11052 10334 11220 10368
rect 11310 10334 11478 10368
rect 11568 10334 11736 10368
rect 11826 10334 11994 10368
rect 12084 10334 12252 10368
rect 12342 10334 12510 10368
rect 12600 10334 12768 10368
rect 10794 9606 10962 9640
rect 11052 9606 11220 9640
rect 11310 9606 11478 9640
rect 11568 9606 11736 9640
rect 11826 9606 11994 9640
rect 12084 9606 12252 9640
rect 12342 9606 12510 9640
rect 12600 9606 12768 9640
rect 13574 11084 13642 11118
rect 13574 10556 13642 10590
rect 14216 11088 14284 11122
rect 14216 9578 14284 9612
<< locali >>
rect 1376 19968 1472 20002
rect 2182 19968 2278 20002
rect 1376 19906 1410 19968
rect 136 18368 232 18402
rect 942 18368 1038 18402
rect 136 18306 170 18368
rect 1004 18306 1038 18368
rect 296 18266 312 18300
rect 350 18266 366 18300
rect 424 18266 440 18300
rect 478 18266 494 18300
rect 552 18266 568 18300
rect 606 18266 622 18300
rect 680 18266 696 18300
rect 734 18266 750 18300
rect 808 18266 824 18300
rect 862 18266 878 18300
rect 250 18207 284 18223
rect 250 16615 284 16631
rect 378 18207 412 18223
rect 378 16615 412 16631
rect 506 18207 540 18223
rect 506 16615 540 16631
rect 634 18207 668 18223
rect 634 16615 668 16631
rect 762 18207 796 18223
rect 762 16615 796 16631
rect 890 18207 924 18223
rect 890 16615 924 16631
rect 296 16538 312 16572
rect 350 16538 366 16572
rect 424 16538 440 16572
rect 478 16538 494 16572
rect 552 16538 568 16572
rect 606 16538 622 16572
rect 680 16538 696 16572
rect 734 16538 750 16572
rect 808 16538 824 16572
rect 862 16538 878 16572
rect 136 16470 170 16532
rect 2244 19906 2278 19968
rect 1536 19866 1552 19900
rect 1590 19866 1606 19900
rect 1664 19866 1680 19900
rect 1718 19866 1734 19900
rect 1792 19866 1808 19900
rect 1846 19866 1862 19900
rect 1920 19866 1936 19900
rect 1974 19866 1990 19900
rect 2048 19866 2064 19900
rect 2102 19866 2118 19900
rect 1490 19807 1524 19823
rect 1490 18215 1524 18231
rect 1618 19807 1652 19823
rect 1618 18215 1652 18231
rect 1746 19807 1780 19823
rect 1746 18215 1780 18231
rect 1874 19807 1908 19823
rect 1874 18215 1908 18231
rect 2002 19807 2036 19823
rect 2002 18215 2036 18231
rect 2130 19807 2164 19823
rect 2130 18215 2164 18231
rect 1536 18138 1552 18172
rect 1590 18138 1606 18172
rect 1664 18138 1680 18172
rect 1718 18138 1734 18172
rect 1792 18138 1808 18172
rect 1846 18138 1862 18172
rect 1920 18138 1936 18172
rect 1974 18138 1990 18172
rect 2048 18138 2064 18172
rect 2102 18138 2118 18172
rect 1376 18070 1410 18132
rect 11885 19375 11981 19409
rect 14209 19375 14305 19409
rect 11885 19313 11919 19375
rect 14271 19313 14305 19375
rect 12091 19241 12107 19275
rect 14083 19241 14099 19275
rect 12023 19213 12057 19229
rect 12023 19129 12057 19145
rect 14133 19213 14167 19229
rect 14133 19129 14167 19145
rect 12091 19083 12107 19117
rect 14083 19083 14099 19117
rect 11885 18983 11919 19045
rect 14271 18983 14305 19045
rect 11885 18949 11981 18983
rect 14209 18949 14305 18983
rect 2244 18070 2278 18132
rect 1376 18036 1472 18070
rect 2182 18036 2278 18070
rect 1004 16470 1038 16532
rect 136 16436 232 16470
rect 942 16436 1038 16470
rect 10890 13926 10986 13960
rect 12902 13926 12998 13960
rect 10890 13864 10924 13926
rect 12964 13864 12998 13926
rect 11070 13788 11086 13822
rect 11254 13788 11270 13822
rect 11328 13788 11344 13822
rect 11512 13788 11528 13822
rect 11586 13788 11602 13822
rect 11770 13788 11786 13822
rect 11844 13788 11860 13822
rect 12028 13788 12044 13822
rect 12102 13788 12118 13822
rect 12286 13788 12302 13822
rect 12360 13788 12376 13822
rect 12544 13788 12560 13822
rect 12618 13788 12634 13822
rect 12802 13788 12818 13822
rect 11024 13738 11058 13754
rect 11024 13146 11058 13162
rect 11282 13738 11316 13754
rect 11282 13146 11316 13162
rect 11540 13738 11574 13754
rect 11540 13146 11574 13162
rect 11798 13738 11832 13754
rect 11798 13146 11832 13162
rect 12056 13738 12090 13754
rect 12056 13146 12090 13162
rect 12314 13738 12348 13754
rect 12314 13146 12348 13162
rect 12572 13738 12606 13754
rect 12572 13146 12606 13162
rect 12830 13738 12864 13754
rect 12830 13146 12864 13162
rect 11070 13078 11086 13112
rect 11254 13078 11270 13112
rect 11328 13078 11344 13112
rect 11512 13078 11528 13112
rect 11586 13078 11602 13112
rect 11770 13078 11786 13112
rect 11844 13078 11860 13112
rect 12028 13078 12044 13112
rect 12102 13078 12118 13112
rect 12286 13078 12302 13112
rect 12360 13078 12376 13112
rect 12544 13078 12560 13112
rect 12618 13078 12634 13112
rect 12802 13078 12818 13112
rect 12964 12974 12998 13036
rect 10890 12940 10986 12974
rect 12902 12940 12998 12974
rect 14020 13126 14116 13160
rect 14384 13126 14480 13160
rect 14020 13064 14054 13126
rect 9308 12722 9404 12756
rect 12868 12722 12964 12756
rect 9308 12660 9342 12722
rect 12930 12660 12964 12722
rect 9488 12584 9504 12618
rect 9672 12584 9688 12618
rect 9746 12584 9762 12618
rect 9930 12584 9946 12618
rect 10004 12584 10020 12618
rect 10188 12584 10204 12618
rect 10262 12584 10278 12618
rect 10446 12584 10462 12618
rect 10520 12584 10536 12618
rect 10704 12584 10720 12618
rect 10778 12584 10794 12618
rect 10962 12584 10978 12618
rect 11036 12584 11052 12618
rect 11220 12584 11236 12618
rect 11294 12584 11310 12618
rect 11478 12584 11494 12618
rect 11552 12584 11568 12618
rect 11736 12584 11752 12618
rect 11810 12584 11826 12618
rect 11994 12584 12010 12618
rect 12068 12584 12084 12618
rect 12252 12584 12268 12618
rect 12326 12584 12342 12618
rect 12510 12584 12526 12618
rect 12584 12584 12600 12618
rect 12768 12584 12784 12618
rect 9442 12525 9476 12541
rect 9442 11933 9476 11949
rect 9700 12525 9734 12541
rect 9700 11933 9734 11949
rect 9958 12525 9992 12541
rect 9958 11933 9992 11949
rect 10216 12525 10250 12541
rect 10216 11933 10250 11949
rect 10474 12525 10508 12541
rect 10474 11933 10508 11949
rect 10732 12525 10766 12541
rect 10732 11933 10766 11949
rect 10990 12525 11024 12541
rect 10990 11933 11024 11949
rect 11248 12525 11282 12541
rect 11248 11933 11282 11949
rect 11506 12525 11540 12541
rect 11506 11933 11540 11949
rect 11764 12525 11798 12541
rect 11764 11933 11798 11949
rect 12022 12525 12056 12541
rect 12022 11933 12056 11949
rect 12280 12525 12314 12541
rect 12280 11933 12314 11949
rect 12538 12525 12572 12541
rect 12538 11933 12572 11949
rect 12796 12525 12830 12541
rect 12796 11933 12830 11949
rect 9488 11856 9504 11890
rect 9672 11856 9688 11890
rect 9746 11856 9762 11890
rect 9930 11856 9946 11890
rect 10004 11856 10020 11890
rect 10188 11856 10204 11890
rect 10262 11856 10278 11890
rect 10446 11856 10462 11890
rect 10520 11856 10536 11890
rect 10704 11856 10720 11890
rect 10778 11856 10794 11890
rect 10962 11856 10978 11890
rect 11036 11856 11052 11890
rect 11220 11856 11236 11890
rect 11294 11856 11310 11890
rect 11478 11856 11494 11890
rect 11552 11856 11568 11890
rect 11736 11856 11752 11890
rect 11810 11856 11826 11890
rect 11994 11856 12010 11890
rect 12068 11856 12084 11890
rect 12252 11856 12268 11890
rect 12326 11856 12342 11890
rect 12510 11856 12526 11890
rect 12584 11856 12600 11890
rect 12768 11856 12784 11890
rect 12930 11752 12964 11814
rect 9308 11718 9404 11752
rect 12868 11718 12964 11752
rect 13378 12142 13474 12176
rect 13742 12142 13838 12176
rect 13378 12080 13412 12142
rect 13804 12080 13838 12142
rect 13558 12004 13574 12038
rect 13642 12004 13658 12038
rect 10598 11602 10694 11636
rect 12868 11602 12964 11636
rect 10598 11540 10632 11602
rect 12930 11540 12964 11602
rect 10778 11464 10794 11498
rect 10962 11464 10978 11498
rect 11036 11464 11052 11498
rect 11220 11464 11236 11498
rect 11294 11464 11310 11498
rect 11478 11464 11494 11498
rect 11552 11464 11568 11498
rect 11736 11464 11752 11498
rect 11810 11464 11826 11498
rect 11994 11464 12010 11498
rect 12068 11464 12084 11498
rect 12252 11464 12268 11498
rect 12326 11464 12342 11498
rect 12510 11464 12526 11498
rect 12584 11464 12600 11498
rect 12768 11464 12784 11498
rect 10732 11405 10766 11421
rect 10732 10813 10766 10829
rect 10990 11405 11024 11421
rect 10990 10813 11024 10829
rect 11248 11405 11282 11421
rect 11248 10813 11282 10829
rect 11506 11405 11540 11421
rect 11506 10813 11540 10829
rect 11764 11405 11798 11421
rect 11764 10813 11798 10829
rect 12022 11405 12056 11421
rect 12022 10813 12056 10829
rect 12280 11405 12314 11421
rect 12280 10813 12314 10829
rect 12538 11405 12572 11421
rect 12538 10813 12572 10829
rect 12796 11405 12830 11421
rect 12796 10813 12830 10829
rect 10778 10736 10794 10770
rect 10962 10736 10978 10770
rect 11036 10736 11052 10770
rect 11220 10736 11236 10770
rect 11294 10736 11310 10770
rect 11478 10736 11494 10770
rect 11552 10736 11568 10770
rect 11736 10736 11752 10770
rect 11810 10736 11826 10770
rect 11994 10736 12010 10770
rect 12068 10736 12084 10770
rect 12252 10736 12268 10770
rect 12326 10736 12342 10770
rect 12510 10736 12526 10770
rect 12584 10736 12600 10770
rect 12768 10736 12784 10770
rect 13512 11945 13546 11961
rect 13512 11553 13546 11569
rect 13670 11945 13704 11961
rect 13670 11553 13704 11569
rect 13558 11476 13574 11510
rect 13642 11476 13658 11510
rect 13378 11372 13412 11434
rect 13804 11372 13838 11434
rect 13378 11338 13474 11372
rect 13742 11338 13838 11372
rect 14446 13064 14480 13126
rect 14200 12988 14216 13022
rect 14284 12988 14300 13022
rect 14154 12938 14188 12954
rect 14154 11546 14188 11562
rect 14312 12938 14346 12954
rect 14312 11546 14346 11562
rect 14200 11478 14216 11512
rect 14284 11478 14300 11512
rect 14020 11374 14054 11436
rect 14020 11340 14116 11374
rect 14384 11340 14480 11374
rect 12930 10632 12964 10694
rect 10598 10598 10694 10632
rect 12868 10598 12964 10632
rect 13378 11222 13474 11256
rect 13742 11222 13838 11256
rect 13378 11160 13412 11222
rect 13804 11160 13838 11222
rect 13558 11084 13574 11118
rect 13642 11084 13658 11118
rect 13512 11025 13546 11041
rect 13512 10633 13546 10649
rect 13670 11025 13704 11041
rect 13670 10633 13704 10649
rect 13558 10556 13574 10590
rect 13642 10556 13658 10590
rect 10598 10472 10694 10506
rect 12868 10472 12964 10506
rect 12930 10410 12964 10472
rect 13378 10452 13412 10514
rect 13804 10452 13838 10514
rect 13378 10418 13474 10452
rect 13742 10418 13838 10452
rect 14020 11226 14116 11260
rect 14384 11226 14480 11260
rect 14020 11164 14054 11226
rect 10778 10334 10794 10368
rect 10962 10334 10978 10368
rect 11036 10334 11052 10368
rect 11220 10334 11236 10368
rect 11294 10334 11310 10368
rect 11478 10334 11494 10368
rect 11552 10334 11568 10368
rect 11736 10334 11752 10368
rect 11810 10334 11826 10368
rect 11994 10334 12010 10368
rect 12068 10334 12084 10368
rect 12252 10334 12268 10368
rect 12326 10334 12342 10368
rect 12510 10334 12526 10368
rect 12584 10334 12600 10368
rect 12768 10334 12784 10368
rect 10732 10275 10766 10291
rect 10732 9683 10766 9699
rect 10990 10275 11024 10291
rect 10990 9683 11024 9699
rect 11248 10275 11282 10291
rect 11248 9683 11282 9699
rect 11506 10275 11540 10291
rect 11506 9683 11540 9699
rect 11764 10275 11798 10291
rect 11764 9683 11798 9699
rect 12022 10275 12056 10291
rect 12022 9683 12056 9699
rect 12280 10275 12314 10291
rect 12280 9683 12314 9699
rect 12538 10275 12572 10291
rect 12538 9683 12572 9699
rect 12796 10275 12830 10291
rect 12796 9683 12830 9699
rect 10778 9606 10794 9640
rect 10962 9606 10978 9640
rect 11036 9606 11052 9640
rect 11220 9606 11236 9640
rect 11294 9606 11310 9640
rect 11478 9606 11494 9640
rect 11552 9606 11568 9640
rect 11736 9606 11752 9640
rect 11810 9606 11826 9640
rect 11994 9606 12010 9640
rect 12068 9606 12084 9640
rect 12252 9606 12268 9640
rect 12326 9606 12342 9640
rect 12510 9606 12526 9640
rect 12584 9606 12600 9640
rect 12768 9606 12784 9640
rect 10598 9502 10632 9564
rect 12930 9502 12964 9564
rect 10598 9468 10694 9502
rect 12868 9468 12964 9502
rect 14200 11088 14216 11122
rect 14284 11088 14300 11122
rect 14154 11038 14188 11054
rect 14154 9646 14188 9662
rect 14312 11038 14346 11054
rect 14312 9646 14346 9662
rect 14200 9578 14216 9612
rect 14284 9578 14300 9612
rect 14020 9474 14054 9536
rect 14446 9474 14480 9536
rect 14020 9440 14116 9474
rect 14384 9440 14480 9474
<< viali >>
rect 1619 19968 2035 20002
rect 379 18368 795 18402
rect 312 18266 350 18300
rect 440 18266 478 18300
rect 568 18266 606 18300
rect 696 18266 734 18300
rect 824 18266 862 18300
rect 250 17560 284 18190
rect 378 16648 412 17278
rect 506 17560 540 18190
rect 634 16648 668 17278
rect 762 17560 796 18190
rect 890 16648 924 17278
rect 312 16538 350 16572
rect 440 16538 478 16572
rect 568 16538 606 16572
rect 696 16538 734 16572
rect 824 16538 862 16572
rect 1552 19866 1590 19900
rect 1680 19866 1718 19900
rect 1808 19866 1846 19900
rect 1936 19866 1974 19900
rect 2064 19866 2102 19900
rect 1490 19160 1524 19790
rect 1618 18248 1652 18878
rect 1746 19160 1780 19790
rect 1874 18248 1908 18878
rect 2002 19160 2036 19790
rect 2130 18248 2164 18878
rect 1552 18138 1590 18172
rect 1680 18138 1718 18172
rect 1808 18138 1846 18172
rect 1936 18138 1974 18172
rect 2064 18138 2102 18172
rect 13671 19241 14066 19275
rect 12023 19145 12057 19213
rect 14133 19145 14167 19213
rect 12124 19083 12519 19117
rect 12919 18949 13271 18983
rect 11086 13788 11254 13822
rect 11344 13788 11512 13822
rect 11602 13788 11770 13822
rect 11860 13788 12028 13822
rect 12118 13788 12286 13822
rect 12376 13788 12544 13822
rect 12634 13788 12802 13822
rect 10890 13036 10924 13450
rect 11024 13491 11058 13721
rect 11282 13179 11316 13409
rect 11540 13491 11574 13721
rect 11798 13179 11832 13409
rect 12056 13491 12090 13721
rect 12314 13179 12348 13409
rect 12572 13491 12606 13721
rect 12830 13179 12864 13409
rect 11086 13078 11254 13112
rect 11344 13078 11512 13112
rect 11602 13078 11770 13112
rect 11860 13078 12028 13112
rect 12118 13078 12286 13112
rect 12376 13078 12544 13112
rect 12634 13078 12802 13112
rect 10890 12974 10924 13036
rect 9504 12584 9672 12618
rect 9762 12584 9930 12618
rect 10020 12584 10188 12618
rect 10278 12584 10446 12618
rect 10536 12584 10704 12618
rect 10794 12584 10962 12618
rect 11052 12584 11220 12618
rect 11310 12584 11478 12618
rect 11568 12584 11736 12618
rect 11826 12584 11994 12618
rect 12084 12584 12252 12618
rect 12342 12584 12510 12618
rect 12600 12584 12768 12618
rect 9308 11814 9342 12237
rect 9442 12278 9476 12508
rect 9700 11966 9734 12196
rect 9958 12278 9992 12508
rect 10216 11966 10250 12196
rect 10474 12278 10508 12508
rect 10732 11966 10766 12196
rect 10990 12278 11024 12508
rect 11248 11966 11282 12196
rect 11506 12278 11540 12508
rect 11764 11966 11798 12196
rect 12022 12278 12056 12508
rect 12280 11966 12314 12196
rect 12538 12278 12572 12508
rect 12796 11966 12830 12196
rect 9504 11856 9672 11890
rect 9762 11856 9930 11890
rect 10020 11856 10188 11890
rect 10278 11856 10446 11890
rect 10536 11856 10704 11890
rect 10794 11856 10962 11890
rect 11052 11856 11220 11890
rect 11310 11856 11478 11890
rect 11568 11856 11736 11890
rect 11826 11856 11994 11890
rect 12084 11856 12252 11890
rect 12342 11856 12510 11890
rect 12600 11856 12768 11890
rect 9308 11752 9342 11814
rect 13574 12004 13642 12038
rect 13378 11699 13412 11815
rect 10794 11464 10962 11498
rect 11052 11464 11220 11498
rect 11310 11464 11478 11498
rect 11568 11464 11736 11498
rect 11826 11464 11994 11498
rect 12084 11464 12252 11498
rect 12342 11464 12510 11498
rect 12600 11464 12768 11498
rect 10598 10694 10632 11117
rect 10732 11158 10766 11388
rect 10990 10846 11024 11076
rect 11248 11158 11282 11388
rect 11506 10846 11540 11076
rect 11764 11158 11798 11388
rect 12022 10846 12056 11076
rect 12280 11158 12314 11388
rect 12538 10846 12572 11076
rect 12796 11158 12830 11388
rect 10794 10736 10962 10770
rect 11052 10736 11220 10770
rect 11310 10736 11478 10770
rect 11568 10736 11736 10770
rect 11826 10736 11994 10770
rect 12084 10736 12252 10770
rect 12342 10736 12510 10770
rect 12600 10736 12768 10770
rect 10598 10632 10632 10694
rect 13512 11569 13546 11945
rect 13670 11569 13704 11945
rect 13574 11476 13642 11510
rect 14216 12988 14284 13022
rect 14154 11579 14188 11992
rect 14312 11579 14346 11992
rect 14216 11478 14284 11512
rect 14446 11436 14480 11900
rect 14446 11374 14480 11436
rect 13574 11084 13642 11118
rect 13378 10779 13412 10895
rect 13512 10649 13546 11025
rect 13670 10649 13704 11025
rect 13574 10556 13642 10590
rect 10598 10410 10632 10472
rect 10598 9987 10632 10410
rect 10794 10334 10962 10368
rect 11052 10334 11220 10368
rect 11310 10334 11478 10368
rect 11568 10334 11736 10368
rect 11826 10334 11994 10368
rect 12084 10334 12252 10368
rect 12342 10334 12510 10368
rect 12600 10334 12768 10368
rect 10732 10028 10766 10258
rect 10990 9716 11024 9946
rect 11248 10028 11282 10258
rect 11506 9716 11540 9946
rect 11764 10028 11798 10258
rect 12022 9716 12056 9946
rect 12280 10028 12314 10258
rect 12538 9716 12572 9946
rect 12796 10028 12830 10258
rect 10794 9606 10962 9640
rect 11052 9606 11220 9640
rect 11310 9606 11478 9640
rect 11568 9606 11736 9640
rect 11826 9606 11994 9640
rect 12084 9606 12252 9640
rect 12342 9606 12510 9640
rect 12600 9606 12768 9640
rect 14446 11164 14480 11226
rect 14216 11088 14284 11122
rect 14154 10608 14188 11021
rect 14312 10608 14346 11021
rect 14446 10700 14480 11164
rect 14216 9578 14284 9612
<< metal1 >>
rect -230 26620 200 26820
rect 0 26600 200 26620
rect 0 26480 40 26600
rect 160 26480 200 26600
rect 0 26440 200 26480
rect 1600 20002 2060 20040
rect 1600 19968 1619 20002
rect 2035 19968 2060 20002
rect 1600 19920 2060 19968
rect 1480 19900 2180 19920
rect 1480 19866 1552 19900
rect 1590 19866 1680 19900
rect 1718 19866 1808 19900
rect 1846 19866 1936 19900
rect 1974 19866 2064 19900
rect 2102 19866 2180 19900
rect 1480 19790 2180 19866
rect 580 19560 740 19580
rect 580 19440 600 19560
rect 720 19440 740 19560
rect 580 18640 740 19440
rect 1480 19160 1490 19790
rect 1524 19160 1746 19790
rect 1780 19160 2002 19790
rect 2036 19740 2180 19790
rect 2036 19720 3300 19740
rect 2036 19560 3120 19720
rect 3280 19560 3300 19720
rect 8900 19720 9330 19740
rect 15000 19720 15430 19740
rect 8900 19700 12370 19720
rect 8640 19680 12370 19700
rect 8640 19580 8660 19680
rect 8780 19580 12370 19680
rect 8640 19560 12370 19580
rect 2036 19540 3300 19560
rect 8900 19540 9330 19560
rect 2036 19160 2180 19540
rect 1480 19140 2180 19160
rect 1612 18878 1658 18890
rect 1612 18640 1618 18878
rect 500 18440 1618 18640
rect 360 18402 820 18440
rect 360 18368 379 18402
rect 795 18368 820 18402
rect 360 18320 820 18368
rect 240 18300 940 18320
rect 240 18266 312 18300
rect 350 18266 440 18300
rect 478 18266 568 18300
rect 606 18266 696 18300
rect 734 18266 824 18300
rect 862 18266 940 18300
rect 240 18190 940 18266
rect 1612 18248 1618 18440
rect 1652 18640 1658 18878
rect 1868 18878 1914 18890
rect 1868 18640 1874 18878
rect 1652 18440 1874 18640
rect 1652 18248 1658 18440
rect 1612 18236 1658 18248
rect 1868 18248 1874 18440
rect 1908 18640 1914 18878
rect 2124 18878 2170 18890
rect 2124 18640 2130 18878
rect 1908 18440 2130 18640
rect 1908 18248 1914 18440
rect 1868 18236 1914 18248
rect 2124 18248 2130 18440
rect 2164 18640 2170 18878
rect 2164 18440 2180 18640
rect 2164 18248 2170 18440
rect 2124 18236 2170 18248
rect 240 17560 250 18190
rect 284 17560 506 18190
rect 540 17560 762 18190
rect 796 17560 940 18190
rect 1540 18172 2120 18180
rect 1540 18138 1552 18172
rect 1590 18138 1680 18172
rect 1718 18138 1808 18172
rect 1846 18138 1936 18172
rect 1974 18138 2064 18172
rect 2102 18138 2120 18172
rect 1540 18120 2120 18138
rect 244 17548 290 17560
rect 500 17548 546 17560
rect 756 17548 802 17560
rect 372 17278 418 17290
rect 372 16940 378 17278
rect 360 16740 378 16940
rect 372 16648 378 16740
rect 412 16940 418 17278
rect 628 17278 674 17290
rect 628 16940 634 17278
rect 412 16740 634 16940
rect 412 16648 418 16740
rect 372 16636 418 16648
rect 628 16648 634 16740
rect 668 16940 674 17278
rect 884 17278 930 17290
rect 884 16940 890 17278
rect 668 16740 890 16940
rect 668 16648 674 16740
rect 628 16636 674 16648
rect 884 16648 890 16740
rect 924 16940 930 17278
rect 924 16740 1180 16940
rect 924 16648 930 16740
rect 884 16636 930 16648
rect 280 16572 880 16580
rect 280 16538 312 16572
rect 350 16538 440 16572
rect 478 16538 568 16572
rect 606 16538 696 16572
rect 734 16538 824 16572
rect 862 16538 880 16572
rect 280 16520 880 16538
rect 980 16380 1180 16740
rect 9150 16650 9310 19540
rect 12017 19213 12063 19225
rect 12017 19145 12023 19213
rect 12057 19145 12063 19213
rect 12017 19133 12063 19145
rect 12220 19123 12370 19560
rect 13790 19700 15430 19720
rect 13790 19580 14560 19700
rect 14680 19580 15430 19700
rect 13790 19560 15430 19580
rect 13790 19281 13940 19560
rect 15000 19540 15430 19560
rect 13659 19275 14078 19281
rect 13659 19241 13671 19275
rect 14066 19241 14078 19275
rect 13659 19235 14078 19241
rect 13790 19230 13940 19235
rect 14130 19225 14700 19230
rect 14127 19213 14700 19225
rect 14127 19145 14133 19213
rect 14167 19145 14700 19213
rect 14127 19133 14700 19145
rect 14130 19130 14700 19133
rect 12112 19117 12531 19123
rect 12112 19083 12124 19117
rect 12519 19083 12531 19117
rect 12112 19077 12531 19083
rect 13030 18989 13160 18990
rect 12907 18983 13283 18989
rect 12907 18949 12919 18983
rect 13271 18949 13283 18983
rect 12907 18943 13283 18949
rect 13030 18910 13160 18943
rect 13030 18820 13050 18910
rect 13140 18820 13160 18910
rect 13030 18800 13160 18820
rect 9150 16530 9170 16650
rect 9290 16530 9310 16650
rect 9150 16510 9310 16530
rect -230 16360 9550 16380
rect -230 16200 2520 16360
rect 2680 16200 9370 16360
rect 9530 16200 9550 16360
rect -230 16180 9550 16200
rect 11074 13822 11266 13828
rect 11074 13788 11086 13822
rect 11254 13788 11266 13822
rect 11074 13782 11266 13788
rect 11332 13822 11524 13828
rect 11332 13788 11344 13822
rect 11512 13788 11524 13822
rect 11332 13782 11524 13788
rect 11590 13822 11782 13828
rect 11590 13788 11602 13822
rect 11770 13788 11782 13822
rect 11590 13782 11782 13788
rect 11848 13822 12040 13828
rect 11848 13788 11860 13822
rect 12028 13788 12040 13822
rect 11848 13782 12040 13788
rect 12106 13822 12298 13828
rect 12106 13788 12118 13822
rect 12286 13788 12298 13822
rect 12106 13782 12298 13788
rect 12364 13822 12556 13828
rect 12364 13788 12376 13822
rect 12544 13788 12556 13822
rect 12364 13782 12556 13788
rect 12622 13822 12814 13828
rect 12622 13788 12634 13822
rect 12802 13788 12814 13822
rect 12622 13782 12814 13788
rect 11018 13721 11064 13733
rect 11018 13680 11024 13721
rect 9150 13530 11024 13680
rect 9150 12470 9310 13530
rect 11018 13491 11024 13530
rect 11058 13680 11064 13721
rect 11534 13721 11580 13733
rect 11534 13680 11540 13721
rect 11058 13530 11540 13680
rect 11058 13491 11064 13530
rect 11018 13479 11064 13491
rect 11534 13491 11540 13530
rect 11574 13680 11580 13721
rect 12050 13721 12096 13733
rect 12050 13680 12056 13721
rect 11574 13530 12056 13680
rect 11574 13491 11580 13530
rect 11534 13479 11580 13491
rect 12050 13491 12056 13530
rect 12090 13680 12096 13721
rect 12566 13721 12612 13733
rect 12566 13680 12572 13721
rect 12090 13530 12572 13680
rect 12090 13491 12096 13530
rect 12050 13479 12096 13491
rect 12566 13491 12572 13530
rect 12606 13680 12612 13721
rect 14540 13710 14700 19130
rect 14520 13680 14720 13710
rect 12606 13660 14720 13680
rect 12606 13550 14360 13660
rect 14460 13550 14720 13660
rect 12606 13530 14720 13550
rect 12606 13491 12612 13530
rect 14520 13510 14720 13530
rect 12566 13479 12612 13491
rect 10884 13450 10930 13462
rect 10884 13370 10890 13450
rect 10880 13220 10890 13370
rect 10884 12974 10890 13220
rect 10924 13370 10930 13450
rect 11276 13409 11322 13421
rect 11276 13370 11282 13409
rect 10924 13220 11282 13370
rect 10924 12974 10930 13220
rect 11276 13179 11282 13220
rect 11316 13370 11322 13409
rect 11792 13409 11838 13421
rect 11792 13370 11798 13409
rect 11316 13220 11798 13370
rect 11316 13179 11322 13220
rect 11276 13167 11322 13179
rect 11792 13179 11798 13220
rect 11832 13370 11838 13409
rect 12308 13409 12354 13421
rect 12308 13370 12314 13409
rect 11832 13220 12314 13370
rect 11832 13179 11838 13220
rect 11792 13167 11838 13179
rect 12308 13179 12314 13220
rect 12348 13370 12354 13409
rect 12824 13409 12870 13421
rect 12824 13370 12830 13409
rect 12348 13220 12830 13370
rect 12348 13179 12354 13220
rect 12308 13167 12354 13179
rect 12824 13179 12830 13220
rect 12864 13370 12870 13409
rect 12864 13350 14700 13370
rect 12864 13240 14560 13350
rect 14680 13240 14700 13350
rect 12864 13220 14700 13240
rect 12864 13179 12870 13220
rect 12824 13167 12870 13179
rect 13460 13120 13470 13130
rect 11070 13112 13470 13120
rect 11070 13078 11086 13112
rect 11254 13078 11344 13112
rect 11512 13078 11602 13112
rect 11770 13078 11860 13112
rect 12028 13078 12118 13112
rect 12286 13078 12376 13112
rect 12544 13078 12634 13112
rect 12802 13078 13470 13112
rect 11070 13050 13470 13078
rect 13460 13040 13470 13050
rect 13560 13040 13570 13130
rect 14204 13022 14296 13028
rect 14204 12988 14216 13022
rect 14284 12988 14296 13022
rect 14204 12982 14296 12988
rect 10884 12962 10930 12974
rect 9492 12618 9684 12624
rect 9492 12584 9504 12618
rect 9672 12584 9684 12618
rect 9492 12578 9684 12584
rect 9750 12618 9942 12624
rect 9750 12584 9762 12618
rect 9930 12584 9942 12618
rect 9750 12578 9942 12584
rect 10008 12618 10200 12624
rect 10008 12584 10020 12618
rect 10188 12584 10200 12618
rect 10008 12578 10200 12584
rect 10266 12618 10458 12624
rect 10266 12584 10278 12618
rect 10446 12584 10458 12618
rect 10266 12578 10458 12584
rect 10524 12618 10716 12624
rect 10524 12584 10536 12618
rect 10704 12584 10716 12618
rect 10524 12578 10716 12584
rect 10782 12618 10974 12624
rect 10782 12584 10794 12618
rect 10962 12584 10974 12618
rect 10782 12578 10974 12584
rect 11040 12618 11232 12624
rect 11040 12584 11052 12618
rect 11220 12584 11232 12618
rect 11040 12578 11232 12584
rect 11298 12618 11490 12624
rect 11298 12584 11310 12618
rect 11478 12584 11490 12618
rect 11298 12578 11490 12584
rect 11556 12618 11748 12624
rect 11556 12584 11568 12618
rect 11736 12584 11748 12618
rect 11556 12578 11748 12584
rect 11814 12618 12006 12624
rect 11814 12584 11826 12618
rect 11994 12584 12006 12618
rect 11814 12578 12006 12584
rect 12072 12618 12264 12624
rect 12072 12584 12084 12618
rect 12252 12584 12264 12618
rect 12072 12578 12264 12584
rect 12330 12618 12522 12624
rect 12330 12584 12342 12618
rect 12510 12584 12522 12618
rect 12330 12578 12522 12584
rect 12588 12618 12780 12624
rect 12588 12584 12600 12618
rect 12768 12584 12780 12618
rect 12588 12578 12780 12584
rect 9436 12508 9482 12520
rect 9436 12470 9442 12508
rect 9150 12320 9442 12470
rect 9436 12278 9442 12320
rect 9476 12470 9482 12508
rect 9952 12508 9998 12520
rect 9952 12470 9958 12508
rect 9476 12320 9958 12470
rect 9476 12278 9482 12320
rect 9436 12266 9482 12278
rect 9952 12278 9958 12320
rect 9992 12470 9998 12508
rect 10468 12508 10514 12520
rect 10468 12470 10474 12508
rect 9992 12320 10474 12470
rect 9992 12278 9998 12320
rect 9952 12266 9998 12278
rect 10468 12278 10474 12320
rect 10508 12470 10514 12508
rect 10984 12508 11030 12520
rect 10984 12470 10990 12508
rect 10508 12320 10990 12470
rect 10508 12278 10514 12320
rect 10468 12266 10514 12278
rect 10984 12278 10990 12320
rect 11024 12470 11030 12508
rect 11500 12508 11546 12520
rect 11500 12470 11506 12508
rect 11024 12320 11506 12470
rect 11024 12278 11030 12320
rect 10984 12266 11030 12278
rect 11500 12278 11506 12320
rect 11540 12470 11546 12508
rect 12016 12508 12062 12520
rect 12016 12470 12022 12508
rect 11540 12320 12022 12470
rect 11540 12278 11546 12320
rect 11500 12266 11546 12278
rect 12016 12278 12022 12320
rect 12056 12470 12062 12508
rect 12532 12508 12578 12520
rect 12532 12470 12538 12508
rect 12056 12320 12538 12470
rect 12056 12278 12062 12320
rect 12016 12266 12062 12278
rect 12532 12278 12538 12320
rect 12572 12470 12578 12508
rect 12572 12320 12580 12470
rect 14520 12390 14720 12410
rect 14970 12390 15400 12410
rect 14520 12360 15400 12390
rect 12572 12278 12578 12320
rect 12532 12266 12578 12278
rect 13560 12260 15400 12360
rect 9302 12237 9348 12249
rect 9302 12150 9308 12237
rect 9150 11752 9308 12150
rect 9342 12150 9348 12237
rect 9694 12196 9740 12208
rect 9694 12150 9700 12196
rect 9342 12000 9700 12150
rect 9342 11752 9348 12000
rect 9694 11966 9700 12000
rect 9734 12150 9740 12196
rect 10210 12196 10256 12208
rect 10210 12150 10216 12196
rect 9734 12000 10216 12150
rect 9734 11966 9740 12000
rect 9694 11954 9740 11966
rect 10210 11966 10216 12000
rect 10250 12150 10256 12196
rect 10726 12196 10772 12208
rect 10726 12150 10732 12196
rect 10250 12000 10732 12150
rect 10250 11966 10256 12000
rect 10210 11954 10256 11966
rect 10726 11966 10732 12000
rect 10766 12150 10772 12196
rect 11242 12196 11288 12208
rect 11242 12150 11248 12196
rect 10766 12000 11248 12150
rect 10766 11966 10772 12000
rect 10726 11954 10772 11966
rect 11242 11966 11248 12000
rect 11282 12150 11288 12196
rect 11758 12196 11804 12208
rect 11758 12150 11764 12196
rect 11282 12000 11764 12150
rect 11282 11966 11288 12000
rect 11242 11954 11288 11966
rect 11758 11966 11764 12000
rect 11798 12150 11804 12196
rect 12274 12196 12320 12208
rect 12274 12150 12280 12196
rect 11798 12000 12280 12150
rect 11798 11966 11804 12000
rect 11758 11954 11804 11966
rect 12274 11966 12280 12000
rect 12314 12150 12320 12196
rect 12790 12196 12836 12208
rect 12790 12150 12796 12196
rect 12314 12000 12796 12150
rect 12314 11966 12320 12000
rect 12274 11954 12320 11966
rect 12790 11966 12796 12000
rect 12830 12150 12836 12196
rect 12830 12000 12840 12150
rect 13560 12038 13660 12260
rect 14520 12230 15400 12260
rect 14520 12210 14720 12230
rect 14970 12210 15400 12230
rect 13560 12004 13574 12038
rect 13642 12004 13660 12038
rect 13560 12000 13660 12004
rect 12830 11966 12836 12000
rect 13562 11998 13654 12000
rect 12790 11954 12836 11966
rect 14148 11992 14194 12004
rect 13506 11945 13552 11957
rect 9490 11890 12790 11910
rect 9490 11856 9504 11890
rect 9672 11856 9762 11890
rect 9930 11856 10020 11890
rect 10188 11856 10278 11890
rect 10446 11856 10536 11890
rect 10704 11856 10794 11890
rect 10962 11856 11052 11890
rect 11220 11856 11310 11890
rect 11478 11856 11568 11890
rect 11736 11856 11826 11890
rect 11994 11856 12084 11890
rect 12252 11856 12342 11890
rect 12510 11856 12600 11890
rect 12768 11856 12790 11890
rect 9490 11820 12790 11856
rect 13506 11830 13512 11945
rect 9150 11740 9348 11752
rect 9150 11490 9310 11740
rect 9150 11370 9170 11490
rect 9290 11370 9310 11490
rect 10340 11530 10430 11820
rect 13280 11815 13512 11830
rect 13280 11699 13378 11815
rect 13412 11699 13512 11815
rect 13280 11680 13512 11699
rect 10340 11520 12790 11530
rect 10340 11450 10350 11520
rect 10420 11498 12790 11520
rect 10420 11464 10794 11498
rect 10962 11464 11052 11498
rect 11220 11464 11310 11498
rect 11478 11464 11568 11498
rect 11736 11464 11826 11498
rect 11994 11464 12084 11498
rect 12252 11464 12342 11498
rect 12510 11464 12600 11498
rect 12768 11464 12790 11498
rect 10420 11450 12790 11464
rect 10340 11440 12790 11450
rect 9150 11070 9310 11370
rect 10726 11388 10772 11400
rect 10726 11158 10732 11388
rect 10766 11350 10772 11388
rect 11242 11388 11288 11400
rect 11242 11350 11248 11388
rect 10766 11200 11248 11350
rect 10766 11158 10772 11200
rect 10726 11146 10772 11158
rect 11242 11158 11248 11200
rect 11282 11350 11288 11388
rect 11758 11388 11804 11400
rect 11758 11350 11764 11388
rect 11282 11200 11764 11350
rect 11282 11158 11288 11200
rect 11242 11146 11288 11158
rect 11758 11158 11764 11200
rect 11798 11350 11804 11388
rect 12274 11388 12320 11400
rect 12274 11350 12280 11388
rect 11798 11200 12280 11350
rect 11798 11158 11804 11200
rect 11758 11146 11804 11158
rect 12274 11158 12280 11200
rect 12314 11350 12320 11388
rect 12790 11388 12836 11400
rect 12790 11350 12796 11388
rect 12314 11200 12796 11350
rect 12314 11158 12320 11200
rect 12274 11146 12320 11158
rect 12790 11158 12796 11200
rect 12830 11350 12836 11388
rect 13280 11350 13360 11680
rect 13506 11569 13512 11680
rect 13546 11569 13552 11945
rect 13506 11557 13552 11569
rect 13664 11945 13710 11957
rect 13664 11569 13670 11945
rect 13704 11830 13710 11945
rect 14148 11830 14154 11992
rect 13704 11810 14154 11830
rect 13704 11700 13900 11810
rect 14010 11700 14154 11810
rect 13704 11680 14154 11700
rect 13704 11569 13710 11680
rect 13664 11557 13710 11569
rect 14148 11579 14154 11680
rect 14188 11579 14194 11992
rect 14148 11567 14194 11579
rect 14306 11992 14352 12004
rect 14306 11579 14312 11992
rect 14346 11830 14352 11992
rect 14440 11900 14486 11912
rect 14440 11830 14446 11900
rect 14346 11680 14446 11830
rect 14346 11579 14352 11680
rect 14306 11567 14352 11579
rect 13562 11510 13654 11516
rect 13562 11476 13574 11510
rect 13642 11476 13654 11510
rect 13562 11470 13654 11476
rect 14200 11512 14300 11520
rect 14200 11478 14216 11512
rect 14284 11478 14300 11512
rect 12830 11200 13360 11350
rect 14200 11330 14300 11478
rect 14440 11374 14446 11680
rect 14480 11830 14486 11900
rect 14480 11810 14700 11830
rect 14480 11700 14560 11810
rect 14680 11700 14700 11810
rect 14480 11680 14700 11700
rect 14480 11374 14486 11680
rect 14540 11400 14700 11680
rect 14770 11810 14930 11830
rect 14770 11700 14790 11810
rect 14910 11700 14930 11810
rect 14440 11362 14486 11374
rect 14520 11380 14720 11400
rect 14770 11380 14930 11700
rect 14970 11380 15170 11400
rect 12830 11158 12836 11200
rect 12790 11146 12836 11158
rect 10592 11117 10638 11129
rect 9130 11040 9330 11070
rect 10592 11040 10598 11117
rect 9130 10890 10598 11040
rect 9130 10870 9330 10890
rect 9150 10220 9310 10870
rect 10592 10632 10598 10890
rect 10632 11040 10638 11117
rect 10984 11076 11030 11088
rect 10984 11040 10990 11076
rect 10632 10890 10990 11040
rect 10632 10632 10638 10890
rect 10984 10846 10990 10890
rect 11024 11040 11030 11076
rect 11500 11076 11546 11088
rect 11500 11040 11506 11076
rect 11024 10890 11506 11040
rect 11024 10846 11030 10890
rect 10984 10834 11030 10846
rect 11500 10846 11506 10890
rect 11540 11040 11546 11076
rect 12016 11076 12062 11088
rect 12016 11040 12022 11076
rect 11540 10890 12022 11040
rect 11540 10846 11546 10890
rect 11500 10834 11546 10846
rect 12016 10846 12022 10890
rect 12056 11040 12062 11076
rect 12532 11076 12578 11088
rect 12532 11040 12538 11076
rect 12056 10890 12538 11040
rect 12056 10846 12062 10890
rect 12016 10834 12062 10846
rect 12532 10846 12538 10890
rect 12572 10846 12578 11076
rect 12532 10834 12578 10846
rect 13280 10910 13360 11200
rect 13900 11270 14300 11330
rect 13562 11118 13654 11124
rect 13562 11084 13574 11118
rect 13642 11084 13654 11118
rect 13562 11078 13654 11084
rect 13506 11025 13552 11037
rect 13506 10910 13512 11025
rect 13280 10895 13512 10910
rect 13280 10779 13378 10895
rect 13412 10779 13512 10895
rect 10782 10770 10974 10776
rect 10782 10736 10794 10770
rect 10962 10736 10974 10770
rect 10782 10730 10974 10736
rect 11040 10770 11232 10776
rect 11040 10736 11052 10770
rect 11220 10736 11232 10770
rect 11040 10730 11232 10736
rect 11298 10770 11490 10776
rect 11298 10736 11310 10770
rect 11478 10736 11490 10770
rect 11298 10730 11490 10736
rect 11556 10770 11748 10776
rect 11556 10736 11568 10770
rect 11736 10736 11748 10770
rect 11556 10730 11748 10736
rect 11814 10770 12006 10776
rect 11814 10736 11826 10770
rect 11994 10736 12006 10770
rect 11814 10730 12006 10736
rect 12072 10770 12264 10776
rect 12072 10736 12084 10770
rect 12252 10736 12264 10770
rect 12072 10730 12264 10736
rect 12330 10770 12522 10776
rect 12330 10736 12342 10770
rect 12510 10736 12522 10770
rect 12330 10730 12522 10736
rect 12588 10770 12780 10776
rect 12588 10736 12600 10770
rect 12768 10736 12780 10770
rect 13280 10760 13512 10779
rect 12588 10730 12780 10736
rect 13506 10649 13512 10760
rect 13546 10649 13552 11025
rect 13506 10637 13552 10649
rect 13664 11025 13710 11037
rect 13664 10649 13670 11025
rect 13704 10910 13710 11025
rect 13900 10910 14000 11270
rect 14200 11122 14300 11270
rect 14200 11088 14216 11122
rect 14284 11088 14300 11122
rect 14200 11080 14300 11088
rect 14440 11226 14486 11238
rect 14148 11021 14194 11033
rect 14148 10910 14154 11021
rect 13704 10760 14154 10910
rect 13704 10649 13710 10760
rect 13664 10637 13710 10649
rect 10592 10620 10638 10632
rect 14148 10608 14154 10760
rect 14188 10608 14194 11021
rect 13560 10590 13660 10600
rect 14148 10596 14194 10608
rect 14306 11021 14352 11033
rect 14306 10608 14312 11021
rect 14346 10910 14352 11021
rect 14440 10910 14446 11226
rect 14346 10760 14446 10910
rect 14346 10608 14352 10760
rect 14440 10700 14446 10760
rect 14480 10910 14486 11226
rect 14520 11220 15170 11380
rect 14520 11200 14720 11220
rect 14970 11200 15170 11220
rect 14540 10910 14700 11200
rect 14480 10760 14700 10910
rect 14480 10700 14486 10760
rect 14440 10688 14486 10700
rect 14306 10596 14352 10608
rect 13560 10556 13574 10590
rect 13642 10556 13660 10590
rect 10592 10472 10638 10484
rect 10592 10220 10598 10472
rect 9150 10070 10598 10220
rect 10592 9987 10598 10070
rect 10632 10220 10638 10472
rect 10782 10368 10974 10374
rect 10782 10334 10794 10368
rect 10962 10334 10974 10368
rect 10782 10328 10974 10334
rect 11040 10368 11232 10374
rect 11040 10334 11052 10368
rect 11220 10334 11232 10368
rect 11040 10328 11232 10334
rect 11298 10368 11490 10374
rect 11298 10334 11310 10368
rect 11478 10334 11490 10368
rect 11298 10328 11490 10334
rect 11556 10368 11748 10374
rect 11556 10334 11568 10368
rect 11736 10334 11748 10368
rect 11556 10328 11748 10334
rect 11814 10368 12006 10374
rect 11814 10334 11826 10368
rect 11994 10334 12006 10368
rect 11814 10328 12006 10334
rect 12072 10368 12264 10374
rect 12072 10334 12084 10368
rect 12252 10334 12264 10368
rect 12072 10328 12264 10334
rect 12330 10368 12522 10374
rect 12330 10334 12342 10368
rect 12510 10334 12522 10368
rect 12330 10328 12522 10334
rect 12588 10368 12780 10374
rect 12588 10334 12600 10368
rect 12768 10334 12780 10368
rect 12588 10328 12780 10334
rect 13560 10340 13660 10556
rect 14540 10520 14700 10540
rect 14540 10410 14560 10520
rect 14680 10410 14700 10520
rect 14540 10390 14700 10410
rect 14520 10340 14720 10390
rect 10726 10258 10772 10270
rect 10726 10220 10732 10258
rect 10632 10070 10732 10220
rect 10632 9987 10638 10070
rect 10726 10028 10732 10070
rect 10766 10220 10772 10258
rect 11242 10258 11288 10270
rect 11242 10220 11248 10258
rect 10766 10070 11248 10220
rect 10766 10028 10772 10070
rect 10726 10016 10772 10028
rect 11242 10028 11248 10070
rect 11282 10220 11288 10258
rect 11758 10258 11804 10270
rect 11758 10220 11764 10258
rect 11282 10070 11764 10220
rect 11282 10028 11288 10070
rect 11242 10016 11288 10028
rect 11758 10028 11764 10070
rect 11798 10220 11804 10258
rect 12274 10258 12320 10270
rect 12274 10220 12280 10258
rect 11798 10070 12280 10220
rect 11798 10028 11804 10070
rect 11758 10016 11804 10028
rect 12274 10028 12280 10070
rect 12314 10220 12320 10258
rect 12790 10258 12836 10270
rect 12790 10220 12796 10258
rect 12314 10070 12796 10220
rect 12314 10028 12320 10070
rect 12274 10016 12320 10028
rect 12790 10028 12796 10070
rect 12830 10028 12836 10258
rect 13560 10240 14720 10340
rect 14520 10190 14720 10240
rect 12790 10016 12836 10028
rect 10592 9975 10638 9987
rect 10984 9946 11030 9958
rect 9130 9910 9330 9940
rect 10984 9910 10990 9946
rect 9130 9880 10990 9910
rect 9130 9790 10340 9880
rect 10430 9790 10990 9880
rect 9130 9760 10990 9790
rect 9130 9740 9330 9760
rect 9150 9490 9310 9740
rect 10340 9670 10430 9760
rect 10984 9716 10990 9760
rect 11024 9910 11030 9946
rect 11500 9946 11546 9958
rect 11500 9910 11506 9946
rect 11024 9760 11506 9910
rect 11024 9716 11030 9760
rect 10984 9704 11030 9716
rect 11500 9716 11506 9760
rect 11540 9910 11546 9946
rect 12016 9946 12062 9958
rect 12016 9910 12022 9946
rect 11540 9760 12022 9910
rect 11540 9716 11546 9760
rect 11500 9704 11546 9716
rect 12016 9716 12022 9760
rect 12056 9910 12062 9946
rect 12532 9946 12578 9958
rect 12532 9910 12538 9946
rect 12056 9760 12538 9910
rect 12056 9716 12062 9760
rect 12016 9704 12062 9716
rect 12532 9716 12538 9760
rect 12572 9910 12578 9946
rect 12572 9760 12580 9910
rect 12572 9716 12578 9760
rect 12532 9704 12578 9716
rect 10340 9640 12790 9670
rect 10340 9606 10794 9640
rect 10962 9606 11052 9640
rect 11220 9606 11310 9640
rect 11478 9606 11568 9640
rect 11736 9606 11826 9640
rect 11994 9606 12084 9640
rect 12252 9606 12342 9640
rect 12510 9606 12600 9640
rect 12768 9606 12790 9640
rect 10340 9580 12790 9606
rect 14204 9612 14296 9618
rect 14204 9578 14216 9612
rect 14284 9578 14296 9612
rect 14204 9572 14296 9578
rect 9130 9290 9330 9490
rect 9150 9140 9310 9290
rect 15200 9140 15400 9160
rect 9150 8980 15400 9140
rect 15200 8960 15400 8980
<< via1 >>
rect 40 26480 160 26600
rect 600 19440 720 19560
rect 3120 19560 3280 19720
rect 8660 19580 8780 19680
rect 14560 19580 14680 19700
rect 13050 18820 13140 18910
rect 9170 16530 9290 16650
rect 2520 16200 2680 16360
rect 9370 16200 9530 16360
rect 14360 13550 14460 13660
rect 14560 13240 14680 13350
rect 13470 13040 13560 13130
rect 9170 11370 9290 11490
rect 10350 11450 10420 11520
rect 13900 11700 14010 11810
rect 14560 11700 14680 11810
rect 14790 11700 14910 11810
rect 14560 10410 14680 10520
rect 10340 9790 10430 9880
<< metal2 >>
rect 40 26600 160 26610
rect 40 26470 160 26480
rect 3120 19720 3280 19730
rect 600 19560 720 19570
rect 14560 19700 14680 19710
rect 8660 19680 8780 19690
rect 8660 19570 8780 19580
rect 14560 19570 14680 19580
rect 3120 19550 3280 19560
rect 600 19430 720 19440
rect 13160 18920 14930 18930
rect 13030 18910 14930 18920
rect 13030 18820 13050 18910
rect 13140 18820 14930 18910
rect 13030 18800 14930 18820
rect 9150 16650 9310 16670
rect 9150 16530 9170 16650
rect 9290 16530 9310 16650
rect 2520 16360 2680 16370
rect 2520 16190 2680 16200
rect 9150 11490 9310 16530
rect 14770 16380 14930 18800
rect 9350 16360 14930 16380
rect 9350 16200 9370 16360
rect 9530 16200 14930 16360
rect 9350 16180 14930 16200
rect 14360 13660 14460 13670
rect 14360 13540 14460 13550
rect 14540 13350 14700 13370
rect 14540 13240 14560 13350
rect 14680 13240 14700 13350
rect 13460 13130 13570 13140
rect 13460 13040 13470 13130
rect 13560 13040 13570 13130
rect 13460 12520 13570 13040
rect 13460 12410 14010 12520
rect 13900 11810 14010 12410
rect 13900 11690 14010 11700
rect 14540 11810 14700 13240
rect 14540 11700 14560 11810
rect 14680 11700 14700 11810
rect 14540 11680 14700 11700
rect 14770 11810 14930 16180
rect 14770 11700 14790 11810
rect 14910 11700 14930 11810
rect 14770 11680 14930 11700
rect 9150 11370 9170 11490
rect 9290 11370 9310 11490
rect 9150 11360 9310 11370
rect 10340 11520 10430 11530
rect 10340 11450 10350 11520
rect 10420 11450 10430 11520
rect 10340 9880 10430 11450
rect 14560 10520 14680 10530
rect 14560 10400 14680 10410
rect 10340 9780 10430 9790
<< via2 >>
rect 40 26480 160 26600
rect 600 19440 720 19560
rect 3120 19560 3280 19720
rect 8660 19580 8780 19680
rect 14560 19580 14680 19700
rect 2520 16200 2680 16360
rect 14360 13550 14460 13660
rect 13470 13040 13560 13130
rect 14560 10410 14680 10520
<< metal3 >>
rect 30 26600 170 26605
rect 30 26480 40 26600
rect 160 26480 170 26600
rect 30 26475 170 26480
rect 100 26252 6399 26280
rect 100 20108 120 26252
rect 184 20108 6399 26252
rect 100 20080 6399 20108
rect 3110 19720 3290 19725
rect 590 19560 730 19565
rect 590 19440 600 19560
rect 720 19440 730 19560
rect 3110 19560 3120 19720
rect 3280 19560 3290 19720
rect 14540 19700 14700 19720
rect 8650 19680 8790 19685
rect 8650 19580 8660 19680
rect 8780 19580 8790 19680
rect 8650 19575 8790 19580
rect 14540 19580 14560 19700
rect 14680 19580 14700 19700
rect 3110 19555 3290 19560
rect 590 19435 730 19440
rect 2700 19422 8999 19450
rect 2700 16385 2720 19422
rect 2690 16365 2720 16385
rect 2510 16360 2720 16365
rect 2510 16200 2520 16360
rect 2680 16200 2720 16360
rect 2510 16195 2720 16200
rect 2690 16175 2720 16195
rect 2700 13278 2720 16175
rect 2784 13278 8999 19422
rect 9560 18802 14459 18830
rect 9560 14058 14375 18802
rect 14439 14058 14459 18802
rect 9560 14030 14459 14058
rect 14350 13660 14470 13665
rect 14350 13550 14360 13660
rect 14460 13550 14470 13660
rect 14350 13545 14470 13550
rect 2700 13250 8999 13278
rect 2700 13122 8999 13150
rect 2700 6978 2720 13122
rect 2784 6978 8999 13122
rect 13460 13130 13570 13135
rect 13460 13040 13470 13130
rect 13560 13040 13570 13130
rect 13460 13035 13570 13040
rect 14540 10520 14700 19580
rect 14540 10410 14560 10520
rect 14680 10410 14700 10520
rect 14540 10390 14700 10410
rect 2700 6950 8999 6978
rect 2700 6822 8999 6850
rect 2700 678 2720 6822
rect 2784 678 8999 6822
rect 2700 650 8999 678
<< via3 >>
rect 40 26480 160 26600
rect 120 20108 184 26252
rect 600 19440 720 19560
rect 3120 19560 3280 19720
rect 8660 19580 8780 19680
rect 2520 16200 2680 16360
rect 2720 13278 2784 19422
rect 14375 14058 14439 18802
rect 14360 13550 14460 13660
rect 2720 6978 2784 13122
rect 13470 13040 13560 13130
rect 2720 678 2784 6822
<< mimcap >>
rect 299 26140 6299 26180
rect 299 20220 339 26140
rect 6259 20220 6299 26140
rect 299 20180 6299 20220
rect 2899 19310 8899 19350
rect 2899 13390 2939 19310
rect 8859 13390 8899 19310
rect 9660 18690 14260 18730
rect 9660 14170 9700 18690
rect 14220 14170 14260 18690
rect 9660 14130 14260 14170
rect 2899 13350 8899 13390
rect 2899 13010 8899 13050
rect 2899 7090 2939 13010
rect 8859 7090 8899 13010
rect 2899 7050 8899 7090
rect 2899 6710 8899 6750
rect 2899 790 2939 6710
rect 8859 790 8899 6710
rect 2899 750 8899 790
<< mimcapcontact >>
rect 339 20220 6259 26140
rect 2939 13390 8859 19310
rect 9700 14170 14220 18690
rect 2939 7090 8859 13010
rect 2939 790 8859 6710
<< metal4 >>
rect 39 26600 161 26601
rect 39 26480 40 26600
rect 160 26480 161 26600
rect 39 26479 161 26480
rect 60 26380 160 26479
rect 60 26280 200 26380
rect 100 26252 200 26280
rect 100 26220 120 26252
rect 104 20108 120 26220
rect 184 20108 200 26252
rect 338 26140 6260 26141
rect 338 20220 339 26140
rect 6259 20220 6260 26140
rect 338 20219 6260 20220
rect 104 20092 200 20108
rect 580 19560 740 20219
rect 580 19440 600 19560
rect 720 19440 740 19560
rect 3100 19720 3300 19740
rect 3100 19560 3120 19720
rect 3280 19560 3300 19720
rect 580 19420 740 19440
rect 2727 19438 2831 19500
rect 2704 19422 2831 19438
rect 2704 16380 2720 19422
rect 2500 16360 2720 16380
rect 2500 16200 2520 16360
rect 2680 16200 2720 16360
rect 2500 16180 2720 16200
rect 2704 13278 2720 16180
rect 2784 13278 2831 19422
rect 3100 19311 3300 19560
rect 8640 19680 8800 19700
rect 8640 19580 8660 19680
rect 8780 19580 8800 19680
rect 5847 19311 5951 19500
rect 8640 19311 8800 19580
rect 2938 19310 8860 19311
rect 2938 13390 2939 19310
rect 8859 13390 8860 19310
rect 14359 18802 14455 18818
rect 9699 18690 14221 18691
rect 9699 14170 9700 18690
rect 14220 14170 14221 18690
rect 9699 14169 14221 14170
rect 2938 13389 8860 13390
rect 2704 13262 2831 13278
rect 2727 13138 2831 13262
rect 2704 13122 2831 13138
rect 2704 6978 2720 13122
rect 2784 6978 2831 13122
rect 5847 13011 5951 13389
rect 13460 13130 13570 14169
rect 14359 14058 14375 18802
rect 14439 14070 14455 18802
rect 14439 14058 14460 14070
rect 14359 14042 14460 14058
rect 14360 13661 14460 14042
rect 14359 13660 14461 13661
rect 14359 13550 14360 13660
rect 14460 13550 14461 13660
rect 14359 13549 14461 13550
rect 13460 13040 13470 13130
rect 13560 13040 13570 13130
rect 13460 13030 13570 13040
rect 2938 13010 8860 13011
rect 2938 7090 2939 13010
rect 8859 7090 8860 13010
rect 2938 7089 8860 7090
rect 2704 6962 2831 6978
rect 2727 6838 2831 6962
rect 2704 6822 2831 6838
rect 2704 678 2720 6822
rect 2784 678 2831 6822
rect 5847 6711 5951 7089
rect 2938 6710 8860 6711
rect 2938 790 2939 6710
rect 8859 790 8860 6710
rect 2938 789 8860 790
rect 2704 662 2831 678
rect 2727 600 2831 662
rect 5847 600 5951 789
<< labels >>
flabel metal1 -230 26620 -30 26820 0 FreeSans 256 0 0 0 top_in
port 0 nsew
flabel metal1 -230 16180 -30 16380 0 FreeSans 256 0 0 0 top_gnd
port 1 nsew
flabel metal1 15230 19540 15430 19740 0 FreeSans 256 0 0 0 top_out
port 4 nsew
flabel metal1 15200 12210 15400 12410 0 FreeSans 256 0 0 0 top_ref
port 3 nsew
flabel metal1 15200 8960 15400 9160 0 FreeSans 256 0 0 0 top_ibias
port 2 nsew
flabel metal1 9130 9290 9330 9490 0 FreeSans 256 0 0 0 x2.ldo_ibias
flabel metal1 9130 19540 9330 19740 0 FreeSans 256 0 0 0 x2.ldo_in
flabel metal1 14970 12210 15170 12410 0 FreeSans 256 0 0 0 x2.ldo_ref
flabel metal1 14970 11200 15170 11400 0 FreeSans 256 0 0 0 x2.ldo_gnd
flabel metal1 15000 19540 15200 19740 0 FreeSans 256 0 0 0 x2.ldo_out
flabel metal1 9130 10870 9330 11070 0 FreeSans 256 0 0 0 x2.x1.VDD
flabel metal1 9130 9740 9330 9940 0 FreeSans 256 0 0 0 x2.x1.Ibias
flabel metal1 14520 11200 14720 11400 0 FreeSans 256 0 0 0 x2.x1.VSS
flabel metal1 14520 13510 14720 13710 0 FreeSans 256 0 0 0 x2.x1.Vout
flabel metal1 14520 12210 14720 12410 0 FreeSans 256 0 0 0 x2.x1.Vip
flabel metal1 14520 10190 14720 10390 0 FreeSans 256 0 0 0 x2.x1.Vin
flabel metal1 0 16180 200 16380 0 FreeSans 256 0 0 0 x1.ground
flabel metal1 0 26620 200 26820 0 FreeSans 256 0 0 0 x1.i
flabel metal1 8900 19540 9100 19740 0 FreeSans 256 0 0 0 x1.o
<< end >>
