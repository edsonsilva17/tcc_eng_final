magic
tech sky130A
magscale 1 2
timestamp 1712932033
<< pwell >>
rect -2569 -1258 2569 1258
<< nnmos >>
rect -2341 -1000 -2241 1000
rect -2183 -1000 -2083 1000
rect -2025 -1000 -1925 1000
rect -1867 -1000 -1767 1000
rect -1709 -1000 -1609 1000
rect -1551 -1000 -1451 1000
rect -1393 -1000 -1293 1000
rect -1235 -1000 -1135 1000
rect -1077 -1000 -977 1000
rect -919 -1000 -819 1000
rect -761 -1000 -661 1000
rect -603 -1000 -503 1000
rect -445 -1000 -345 1000
rect -287 -1000 -187 1000
rect -129 -1000 -29 1000
rect 29 -1000 129 1000
rect 187 -1000 287 1000
rect 345 -1000 445 1000
rect 503 -1000 603 1000
rect 661 -1000 761 1000
rect 819 -1000 919 1000
rect 977 -1000 1077 1000
rect 1135 -1000 1235 1000
rect 1293 -1000 1393 1000
rect 1451 -1000 1551 1000
rect 1609 -1000 1709 1000
rect 1767 -1000 1867 1000
rect 1925 -1000 2025 1000
rect 2083 -1000 2183 1000
rect 2241 -1000 2341 1000
<< mvndiff >>
rect -2399 988 -2341 1000
rect -2399 -988 -2387 988
rect -2353 -988 -2341 988
rect -2399 -1000 -2341 -988
rect -2241 988 -2183 1000
rect -2241 -988 -2229 988
rect -2195 -988 -2183 988
rect -2241 -1000 -2183 -988
rect -2083 988 -2025 1000
rect -2083 -988 -2071 988
rect -2037 -988 -2025 988
rect -2083 -1000 -2025 -988
rect -1925 988 -1867 1000
rect -1925 -988 -1913 988
rect -1879 -988 -1867 988
rect -1925 -1000 -1867 -988
rect -1767 988 -1709 1000
rect -1767 -988 -1755 988
rect -1721 -988 -1709 988
rect -1767 -1000 -1709 -988
rect -1609 988 -1551 1000
rect -1609 -988 -1597 988
rect -1563 -988 -1551 988
rect -1609 -1000 -1551 -988
rect -1451 988 -1393 1000
rect -1451 -988 -1439 988
rect -1405 -988 -1393 988
rect -1451 -1000 -1393 -988
rect -1293 988 -1235 1000
rect -1293 -988 -1281 988
rect -1247 -988 -1235 988
rect -1293 -1000 -1235 -988
rect -1135 988 -1077 1000
rect -1135 -988 -1123 988
rect -1089 -988 -1077 988
rect -1135 -1000 -1077 -988
rect -977 988 -919 1000
rect -977 -988 -965 988
rect -931 -988 -919 988
rect -977 -1000 -919 -988
rect -819 988 -761 1000
rect -819 -988 -807 988
rect -773 -988 -761 988
rect -819 -1000 -761 -988
rect -661 988 -603 1000
rect -661 -988 -649 988
rect -615 -988 -603 988
rect -661 -1000 -603 -988
rect -503 988 -445 1000
rect -503 -988 -491 988
rect -457 -988 -445 988
rect -503 -1000 -445 -988
rect -345 988 -287 1000
rect -345 -988 -333 988
rect -299 -988 -287 988
rect -345 -1000 -287 -988
rect -187 988 -129 1000
rect -187 -988 -175 988
rect -141 -988 -129 988
rect -187 -1000 -129 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 129 988 187 1000
rect 129 -988 141 988
rect 175 -988 187 988
rect 129 -1000 187 -988
rect 287 988 345 1000
rect 287 -988 299 988
rect 333 -988 345 988
rect 287 -1000 345 -988
rect 445 988 503 1000
rect 445 -988 457 988
rect 491 -988 503 988
rect 445 -1000 503 -988
rect 603 988 661 1000
rect 603 -988 615 988
rect 649 -988 661 988
rect 603 -1000 661 -988
rect 761 988 819 1000
rect 761 -988 773 988
rect 807 -988 819 988
rect 761 -1000 819 -988
rect 919 988 977 1000
rect 919 -988 931 988
rect 965 -988 977 988
rect 919 -1000 977 -988
rect 1077 988 1135 1000
rect 1077 -988 1089 988
rect 1123 -988 1135 988
rect 1077 -1000 1135 -988
rect 1235 988 1293 1000
rect 1235 -988 1247 988
rect 1281 -988 1293 988
rect 1235 -1000 1293 -988
rect 1393 988 1451 1000
rect 1393 -988 1405 988
rect 1439 -988 1451 988
rect 1393 -1000 1451 -988
rect 1551 988 1609 1000
rect 1551 -988 1563 988
rect 1597 -988 1609 988
rect 1551 -1000 1609 -988
rect 1709 988 1767 1000
rect 1709 -988 1721 988
rect 1755 -988 1767 988
rect 1709 -1000 1767 -988
rect 1867 988 1925 1000
rect 1867 -988 1879 988
rect 1913 -988 1925 988
rect 1867 -1000 1925 -988
rect 2025 988 2083 1000
rect 2025 -988 2037 988
rect 2071 -988 2083 988
rect 2025 -1000 2083 -988
rect 2183 988 2241 1000
rect 2183 -988 2195 988
rect 2229 -988 2241 988
rect 2183 -1000 2241 -988
rect 2341 988 2399 1000
rect 2341 -988 2353 988
rect 2387 -988 2399 988
rect 2341 -1000 2399 -988
<< mvndiffc >>
rect -2387 -988 -2353 988
rect -2229 -988 -2195 988
rect -2071 -988 -2037 988
rect -1913 -988 -1879 988
rect -1755 -988 -1721 988
rect -1597 -988 -1563 988
rect -1439 -988 -1405 988
rect -1281 -988 -1247 988
rect -1123 -988 -1089 988
rect -965 -988 -931 988
rect -807 -988 -773 988
rect -649 -988 -615 988
rect -491 -988 -457 988
rect -333 -988 -299 988
rect -175 -988 -141 988
rect -17 -988 17 988
rect 141 -988 175 988
rect 299 -988 333 988
rect 457 -988 491 988
rect 615 -988 649 988
rect 773 -988 807 988
rect 931 -988 965 988
rect 1089 -988 1123 988
rect 1247 -988 1281 988
rect 1405 -988 1439 988
rect 1563 -988 1597 988
rect 1721 -988 1755 988
rect 1879 -988 1913 988
rect 2037 -988 2071 988
rect 2195 -988 2229 988
rect 2353 -988 2387 988
<< mvpsubdiff >>
rect -2533 1210 2533 1222
rect -2533 1176 -2425 1210
rect 2425 1176 2533 1210
rect -2533 1164 2533 1176
rect -2533 1114 -2475 1164
rect -2533 -1114 -2521 1114
rect -2487 -1114 -2475 1114
rect 2475 1114 2533 1164
rect -2533 -1164 -2475 -1114
rect 2475 -1114 2487 1114
rect 2521 -1114 2533 1114
rect 2475 -1164 2533 -1114
rect -2533 -1176 2533 -1164
rect -2533 -1210 -2425 -1176
rect 2425 -1210 2533 -1176
rect -2533 -1222 2533 -1210
<< mvpsubdiffcont >>
rect -2425 1176 2425 1210
rect -2521 -1114 -2487 1114
rect 2487 -1114 2521 1114
rect -2425 -1210 2425 -1176
<< poly >>
rect -2341 1072 -2241 1088
rect -2341 1038 -2325 1072
rect -2257 1038 -2241 1072
rect -2341 1000 -2241 1038
rect -2183 1072 -2083 1088
rect -2183 1038 -2167 1072
rect -2099 1038 -2083 1072
rect -2183 1000 -2083 1038
rect -2025 1072 -1925 1088
rect -2025 1038 -2009 1072
rect -1941 1038 -1925 1072
rect -2025 1000 -1925 1038
rect -1867 1072 -1767 1088
rect -1867 1038 -1851 1072
rect -1783 1038 -1767 1072
rect -1867 1000 -1767 1038
rect -1709 1072 -1609 1088
rect -1709 1038 -1693 1072
rect -1625 1038 -1609 1072
rect -1709 1000 -1609 1038
rect -1551 1072 -1451 1088
rect -1551 1038 -1535 1072
rect -1467 1038 -1451 1072
rect -1551 1000 -1451 1038
rect -1393 1072 -1293 1088
rect -1393 1038 -1377 1072
rect -1309 1038 -1293 1072
rect -1393 1000 -1293 1038
rect -1235 1072 -1135 1088
rect -1235 1038 -1219 1072
rect -1151 1038 -1135 1072
rect -1235 1000 -1135 1038
rect -1077 1072 -977 1088
rect -1077 1038 -1061 1072
rect -993 1038 -977 1072
rect -1077 1000 -977 1038
rect -919 1072 -819 1088
rect -919 1038 -903 1072
rect -835 1038 -819 1072
rect -919 1000 -819 1038
rect -761 1072 -661 1088
rect -761 1038 -745 1072
rect -677 1038 -661 1072
rect -761 1000 -661 1038
rect -603 1072 -503 1088
rect -603 1038 -587 1072
rect -519 1038 -503 1072
rect -603 1000 -503 1038
rect -445 1072 -345 1088
rect -445 1038 -429 1072
rect -361 1038 -345 1072
rect -445 1000 -345 1038
rect -287 1072 -187 1088
rect -287 1038 -271 1072
rect -203 1038 -187 1072
rect -287 1000 -187 1038
rect -129 1072 -29 1088
rect -129 1038 -113 1072
rect -45 1038 -29 1072
rect -129 1000 -29 1038
rect 29 1072 129 1088
rect 29 1038 45 1072
rect 113 1038 129 1072
rect 29 1000 129 1038
rect 187 1072 287 1088
rect 187 1038 203 1072
rect 271 1038 287 1072
rect 187 1000 287 1038
rect 345 1072 445 1088
rect 345 1038 361 1072
rect 429 1038 445 1072
rect 345 1000 445 1038
rect 503 1072 603 1088
rect 503 1038 519 1072
rect 587 1038 603 1072
rect 503 1000 603 1038
rect 661 1072 761 1088
rect 661 1038 677 1072
rect 745 1038 761 1072
rect 661 1000 761 1038
rect 819 1072 919 1088
rect 819 1038 835 1072
rect 903 1038 919 1072
rect 819 1000 919 1038
rect 977 1072 1077 1088
rect 977 1038 993 1072
rect 1061 1038 1077 1072
rect 977 1000 1077 1038
rect 1135 1072 1235 1088
rect 1135 1038 1151 1072
rect 1219 1038 1235 1072
rect 1135 1000 1235 1038
rect 1293 1072 1393 1088
rect 1293 1038 1309 1072
rect 1377 1038 1393 1072
rect 1293 1000 1393 1038
rect 1451 1072 1551 1088
rect 1451 1038 1467 1072
rect 1535 1038 1551 1072
rect 1451 1000 1551 1038
rect 1609 1072 1709 1088
rect 1609 1038 1625 1072
rect 1693 1038 1709 1072
rect 1609 1000 1709 1038
rect 1767 1072 1867 1088
rect 1767 1038 1783 1072
rect 1851 1038 1867 1072
rect 1767 1000 1867 1038
rect 1925 1072 2025 1088
rect 1925 1038 1941 1072
rect 2009 1038 2025 1072
rect 1925 1000 2025 1038
rect 2083 1072 2183 1088
rect 2083 1038 2099 1072
rect 2167 1038 2183 1072
rect 2083 1000 2183 1038
rect 2241 1072 2341 1088
rect 2241 1038 2257 1072
rect 2325 1038 2341 1072
rect 2241 1000 2341 1038
rect -2341 -1038 -2241 -1000
rect -2341 -1072 -2325 -1038
rect -2257 -1072 -2241 -1038
rect -2341 -1088 -2241 -1072
rect -2183 -1038 -2083 -1000
rect -2183 -1072 -2167 -1038
rect -2099 -1072 -2083 -1038
rect -2183 -1088 -2083 -1072
rect -2025 -1038 -1925 -1000
rect -2025 -1072 -2009 -1038
rect -1941 -1072 -1925 -1038
rect -2025 -1088 -1925 -1072
rect -1867 -1038 -1767 -1000
rect -1867 -1072 -1851 -1038
rect -1783 -1072 -1767 -1038
rect -1867 -1088 -1767 -1072
rect -1709 -1038 -1609 -1000
rect -1709 -1072 -1693 -1038
rect -1625 -1072 -1609 -1038
rect -1709 -1088 -1609 -1072
rect -1551 -1038 -1451 -1000
rect -1551 -1072 -1535 -1038
rect -1467 -1072 -1451 -1038
rect -1551 -1088 -1451 -1072
rect -1393 -1038 -1293 -1000
rect -1393 -1072 -1377 -1038
rect -1309 -1072 -1293 -1038
rect -1393 -1088 -1293 -1072
rect -1235 -1038 -1135 -1000
rect -1235 -1072 -1219 -1038
rect -1151 -1072 -1135 -1038
rect -1235 -1088 -1135 -1072
rect -1077 -1038 -977 -1000
rect -1077 -1072 -1061 -1038
rect -993 -1072 -977 -1038
rect -1077 -1088 -977 -1072
rect -919 -1038 -819 -1000
rect -919 -1072 -903 -1038
rect -835 -1072 -819 -1038
rect -919 -1088 -819 -1072
rect -761 -1038 -661 -1000
rect -761 -1072 -745 -1038
rect -677 -1072 -661 -1038
rect -761 -1088 -661 -1072
rect -603 -1038 -503 -1000
rect -603 -1072 -587 -1038
rect -519 -1072 -503 -1038
rect -603 -1088 -503 -1072
rect -445 -1038 -345 -1000
rect -445 -1072 -429 -1038
rect -361 -1072 -345 -1038
rect -445 -1088 -345 -1072
rect -287 -1038 -187 -1000
rect -287 -1072 -271 -1038
rect -203 -1072 -187 -1038
rect -287 -1088 -187 -1072
rect -129 -1038 -29 -1000
rect -129 -1072 -113 -1038
rect -45 -1072 -29 -1038
rect -129 -1088 -29 -1072
rect 29 -1038 129 -1000
rect 29 -1072 45 -1038
rect 113 -1072 129 -1038
rect 29 -1088 129 -1072
rect 187 -1038 287 -1000
rect 187 -1072 203 -1038
rect 271 -1072 287 -1038
rect 187 -1088 287 -1072
rect 345 -1038 445 -1000
rect 345 -1072 361 -1038
rect 429 -1072 445 -1038
rect 345 -1088 445 -1072
rect 503 -1038 603 -1000
rect 503 -1072 519 -1038
rect 587 -1072 603 -1038
rect 503 -1088 603 -1072
rect 661 -1038 761 -1000
rect 661 -1072 677 -1038
rect 745 -1072 761 -1038
rect 661 -1088 761 -1072
rect 819 -1038 919 -1000
rect 819 -1072 835 -1038
rect 903 -1072 919 -1038
rect 819 -1088 919 -1072
rect 977 -1038 1077 -1000
rect 977 -1072 993 -1038
rect 1061 -1072 1077 -1038
rect 977 -1088 1077 -1072
rect 1135 -1038 1235 -1000
rect 1135 -1072 1151 -1038
rect 1219 -1072 1235 -1038
rect 1135 -1088 1235 -1072
rect 1293 -1038 1393 -1000
rect 1293 -1072 1309 -1038
rect 1377 -1072 1393 -1038
rect 1293 -1088 1393 -1072
rect 1451 -1038 1551 -1000
rect 1451 -1072 1467 -1038
rect 1535 -1072 1551 -1038
rect 1451 -1088 1551 -1072
rect 1609 -1038 1709 -1000
rect 1609 -1072 1625 -1038
rect 1693 -1072 1709 -1038
rect 1609 -1088 1709 -1072
rect 1767 -1038 1867 -1000
rect 1767 -1072 1783 -1038
rect 1851 -1072 1867 -1038
rect 1767 -1088 1867 -1072
rect 1925 -1038 2025 -1000
rect 1925 -1072 1941 -1038
rect 2009 -1072 2025 -1038
rect 1925 -1088 2025 -1072
rect 2083 -1038 2183 -1000
rect 2083 -1072 2099 -1038
rect 2167 -1072 2183 -1038
rect 2083 -1088 2183 -1072
rect 2241 -1038 2341 -1000
rect 2241 -1072 2257 -1038
rect 2325 -1072 2341 -1038
rect 2241 -1088 2341 -1072
<< polycont >>
rect -2325 1038 -2257 1072
rect -2167 1038 -2099 1072
rect -2009 1038 -1941 1072
rect -1851 1038 -1783 1072
rect -1693 1038 -1625 1072
rect -1535 1038 -1467 1072
rect -1377 1038 -1309 1072
rect -1219 1038 -1151 1072
rect -1061 1038 -993 1072
rect -903 1038 -835 1072
rect -745 1038 -677 1072
rect -587 1038 -519 1072
rect -429 1038 -361 1072
rect -271 1038 -203 1072
rect -113 1038 -45 1072
rect 45 1038 113 1072
rect 203 1038 271 1072
rect 361 1038 429 1072
rect 519 1038 587 1072
rect 677 1038 745 1072
rect 835 1038 903 1072
rect 993 1038 1061 1072
rect 1151 1038 1219 1072
rect 1309 1038 1377 1072
rect 1467 1038 1535 1072
rect 1625 1038 1693 1072
rect 1783 1038 1851 1072
rect 1941 1038 2009 1072
rect 2099 1038 2167 1072
rect 2257 1038 2325 1072
rect -2325 -1072 -2257 -1038
rect -2167 -1072 -2099 -1038
rect -2009 -1072 -1941 -1038
rect -1851 -1072 -1783 -1038
rect -1693 -1072 -1625 -1038
rect -1535 -1072 -1467 -1038
rect -1377 -1072 -1309 -1038
rect -1219 -1072 -1151 -1038
rect -1061 -1072 -993 -1038
rect -903 -1072 -835 -1038
rect -745 -1072 -677 -1038
rect -587 -1072 -519 -1038
rect -429 -1072 -361 -1038
rect -271 -1072 -203 -1038
rect -113 -1072 -45 -1038
rect 45 -1072 113 -1038
rect 203 -1072 271 -1038
rect 361 -1072 429 -1038
rect 519 -1072 587 -1038
rect 677 -1072 745 -1038
rect 835 -1072 903 -1038
rect 993 -1072 1061 -1038
rect 1151 -1072 1219 -1038
rect 1309 -1072 1377 -1038
rect 1467 -1072 1535 -1038
rect 1625 -1072 1693 -1038
rect 1783 -1072 1851 -1038
rect 1941 -1072 2009 -1038
rect 2099 -1072 2167 -1038
rect 2257 -1072 2325 -1038
<< locali >>
rect -2521 1176 -2425 1210
rect 2425 1176 2521 1210
rect -2521 1114 -2487 1176
rect 2487 1114 2521 1176
rect -2341 1038 -2325 1072
rect -2257 1038 -2241 1072
rect -2183 1038 -2167 1072
rect -2099 1038 -2083 1072
rect -2025 1038 -2009 1072
rect -1941 1038 -1925 1072
rect -1867 1038 -1851 1072
rect -1783 1038 -1767 1072
rect -1709 1038 -1693 1072
rect -1625 1038 -1609 1072
rect -1551 1038 -1535 1072
rect -1467 1038 -1451 1072
rect -1393 1038 -1377 1072
rect -1309 1038 -1293 1072
rect -1235 1038 -1219 1072
rect -1151 1038 -1135 1072
rect -1077 1038 -1061 1072
rect -993 1038 -977 1072
rect -919 1038 -903 1072
rect -835 1038 -819 1072
rect -761 1038 -745 1072
rect -677 1038 -661 1072
rect -603 1038 -587 1072
rect -519 1038 -503 1072
rect -445 1038 -429 1072
rect -361 1038 -345 1072
rect -287 1038 -271 1072
rect -203 1038 -187 1072
rect -129 1038 -113 1072
rect -45 1038 -29 1072
rect 29 1038 45 1072
rect 113 1038 129 1072
rect 187 1038 203 1072
rect 271 1038 287 1072
rect 345 1038 361 1072
rect 429 1038 445 1072
rect 503 1038 519 1072
rect 587 1038 603 1072
rect 661 1038 677 1072
rect 745 1038 761 1072
rect 819 1038 835 1072
rect 903 1038 919 1072
rect 977 1038 993 1072
rect 1061 1038 1077 1072
rect 1135 1038 1151 1072
rect 1219 1038 1235 1072
rect 1293 1038 1309 1072
rect 1377 1038 1393 1072
rect 1451 1038 1467 1072
rect 1535 1038 1551 1072
rect 1609 1038 1625 1072
rect 1693 1038 1709 1072
rect 1767 1038 1783 1072
rect 1851 1038 1867 1072
rect 1925 1038 1941 1072
rect 2009 1038 2025 1072
rect 2083 1038 2099 1072
rect 2167 1038 2183 1072
rect 2241 1038 2257 1072
rect 2325 1038 2341 1072
rect -2387 988 -2353 1004
rect -2387 -1004 -2353 -988
rect -2229 988 -2195 1004
rect -2229 -1004 -2195 -988
rect -2071 988 -2037 1004
rect -2071 -1004 -2037 -988
rect -1913 988 -1879 1004
rect -1913 -1004 -1879 -988
rect -1755 988 -1721 1004
rect -1755 -1004 -1721 -988
rect -1597 988 -1563 1004
rect -1597 -1004 -1563 -988
rect -1439 988 -1405 1004
rect -1439 -1004 -1405 -988
rect -1281 988 -1247 1004
rect -1281 -1004 -1247 -988
rect -1123 988 -1089 1004
rect -1123 -1004 -1089 -988
rect -965 988 -931 1004
rect -965 -1004 -931 -988
rect -807 988 -773 1004
rect -807 -1004 -773 -988
rect -649 988 -615 1004
rect -649 -1004 -615 -988
rect -491 988 -457 1004
rect -491 -1004 -457 -988
rect -333 988 -299 1004
rect -333 -1004 -299 -988
rect -175 988 -141 1004
rect -175 -1004 -141 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 141 988 175 1004
rect 141 -1004 175 -988
rect 299 988 333 1004
rect 299 -1004 333 -988
rect 457 988 491 1004
rect 457 -1004 491 -988
rect 615 988 649 1004
rect 615 -1004 649 -988
rect 773 988 807 1004
rect 773 -1004 807 -988
rect 931 988 965 1004
rect 931 -1004 965 -988
rect 1089 988 1123 1004
rect 1089 -1004 1123 -988
rect 1247 988 1281 1004
rect 1247 -1004 1281 -988
rect 1405 988 1439 1004
rect 1405 -1004 1439 -988
rect 1563 988 1597 1004
rect 1563 -1004 1597 -988
rect 1721 988 1755 1004
rect 1721 -1004 1755 -988
rect 1879 988 1913 1004
rect 1879 -1004 1913 -988
rect 2037 988 2071 1004
rect 2037 -1004 2071 -988
rect 2195 988 2229 1004
rect 2195 -1004 2229 -988
rect 2353 988 2387 1004
rect 2353 -1004 2387 -988
rect -2341 -1072 -2325 -1038
rect -2257 -1072 -2241 -1038
rect -2183 -1072 -2167 -1038
rect -2099 -1072 -2083 -1038
rect -2025 -1072 -2009 -1038
rect -1941 -1072 -1925 -1038
rect -1867 -1072 -1851 -1038
rect -1783 -1072 -1767 -1038
rect -1709 -1072 -1693 -1038
rect -1625 -1072 -1609 -1038
rect -1551 -1072 -1535 -1038
rect -1467 -1072 -1451 -1038
rect -1393 -1072 -1377 -1038
rect -1309 -1072 -1293 -1038
rect -1235 -1072 -1219 -1038
rect -1151 -1072 -1135 -1038
rect -1077 -1072 -1061 -1038
rect -993 -1072 -977 -1038
rect -919 -1072 -903 -1038
rect -835 -1072 -819 -1038
rect -761 -1072 -745 -1038
rect -677 -1072 -661 -1038
rect -603 -1072 -587 -1038
rect -519 -1072 -503 -1038
rect -445 -1072 -429 -1038
rect -361 -1072 -345 -1038
rect -287 -1072 -271 -1038
rect -203 -1072 -187 -1038
rect -129 -1072 -113 -1038
rect -45 -1072 -29 -1038
rect 29 -1072 45 -1038
rect 113 -1072 129 -1038
rect 187 -1072 203 -1038
rect 271 -1072 287 -1038
rect 345 -1072 361 -1038
rect 429 -1072 445 -1038
rect 503 -1072 519 -1038
rect 587 -1072 603 -1038
rect 661 -1072 677 -1038
rect 745 -1072 761 -1038
rect 819 -1072 835 -1038
rect 903 -1072 919 -1038
rect 977 -1072 993 -1038
rect 1061 -1072 1077 -1038
rect 1135 -1072 1151 -1038
rect 1219 -1072 1235 -1038
rect 1293 -1072 1309 -1038
rect 1377 -1072 1393 -1038
rect 1451 -1072 1467 -1038
rect 1535 -1072 1551 -1038
rect 1609 -1072 1625 -1038
rect 1693 -1072 1709 -1038
rect 1767 -1072 1783 -1038
rect 1851 -1072 1867 -1038
rect 1925 -1072 1941 -1038
rect 2009 -1072 2025 -1038
rect 2083 -1072 2099 -1038
rect 2167 -1072 2183 -1038
rect 2241 -1072 2257 -1038
rect 2325 -1072 2341 -1038
rect -2521 -1176 -2487 -1114
rect 2487 -1176 2521 -1114
rect -2521 -1210 -2425 -1176
rect 2425 -1210 2521 -1176
<< viali >>
rect -2325 1038 -2257 1072
rect -2167 1038 -2099 1072
rect -2009 1038 -1941 1072
rect -1851 1038 -1783 1072
rect -1693 1038 -1625 1072
rect -1535 1038 -1467 1072
rect -1377 1038 -1309 1072
rect -1219 1038 -1151 1072
rect -1061 1038 -993 1072
rect -903 1038 -835 1072
rect -745 1038 -677 1072
rect -587 1038 -519 1072
rect -429 1038 -361 1072
rect -271 1038 -203 1072
rect -113 1038 -45 1072
rect 45 1038 113 1072
rect 203 1038 271 1072
rect 361 1038 429 1072
rect 519 1038 587 1072
rect 677 1038 745 1072
rect 835 1038 903 1072
rect 993 1038 1061 1072
rect 1151 1038 1219 1072
rect 1309 1038 1377 1072
rect 1467 1038 1535 1072
rect 1625 1038 1693 1072
rect 1783 1038 1851 1072
rect 1941 1038 2009 1072
rect 2099 1038 2167 1072
rect 2257 1038 2325 1072
rect -2387 -971 -2353 -181
rect -2229 181 -2195 971
rect -2071 -971 -2037 -181
rect -1913 181 -1879 971
rect -1755 -971 -1721 -181
rect -1597 181 -1563 971
rect -1439 -971 -1405 -181
rect -1281 181 -1247 971
rect -1123 -971 -1089 -181
rect -965 181 -931 971
rect -807 -971 -773 -181
rect -649 181 -615 971
rect -491 -971 -457 -181
rect -333 181 -299 971
rect -175 -971 -141 -181
rect -17 181 17 971
rect 141 -971 175 -181
rect 299 181 333 971
rect 457 -971 491 -181
rect 615 181 649 971
rect 773 -971 807 -181
rect 931 181 965 971
rect 1089 -971 1123 -181
rect 1247 181 1281 971
rect 1405 -971 1439 -181
rect 1563 181 1597 971
rect 1721 -971 1755 -181
rect 1879 181 1913 971
rect 2037 -971 2071 -181
rect 2195 181 2229 971
rect 2353 -971 2387 -181
rect -2325 -1072 -2257 -1038
rect -2167 -1072 -2099 -1038
rect -2009 -1072 -1941 -1038
rect -1851 -1072 -1783 -1038
rect -1693 -1072 -1625 -1038
rect -1535 -1072 -1467 -1038
rect -1377 -1072 -1309 -1038
rect -1219 -1072 -1151 -1038
rect -1061 -1072 -993 -1038
rect -903 -1072 -835 -1038
rect -745 -1072 -677 -1038
rect -587 -1072 -519 -1038
rect -429 -1072 -361 -1038
rect -271 -1072 -203 -1038
rect -113 -1072 -45 -1038
rect 45 -1072 113 -1038
rect 203 -1072 271 -1038
rect 361 -1072 429 -1038
rect 519 -1072 587 -1038
rect 677 -1072 745 -1038
rect 835 -1072 903 -1038
rect 993 -1072 1061 -1038
rect 1151 -1072 1219 -1038
rect 1309 -1072 1377 -1038
rect 1467 -1072 1535 -1038
rect 1625 -1072 1693 -1038
rect 1783 -1072 1851 -1038
rect 1941 -1072 2009 -1038
rect 2099 -1072 2167 -1038
rect 2257 -1072 2325 -1038
rect -124 -1210 124 -1176
<< metal1 >>
rect -2337 1072 -2245 1078
rect -2337 1038 -2325 1072
rect -2257 1038 -2245 1072
rect -2337 1032 -2245 1038
rect -2179 1072 -2087 1078
rect -2179 1038 -2167 1072
rect -2099 1038 -2087 1072
rect -2179 1032 -2087 1038
rect -2021 1072 -1929 1078
rect -2021 1038 -2009 1072
rect -1941 1038 -1929 1072
rect -2021 1032 -1929 1038
rect -1863 1072 -1771 1078
rect -1863 1038 -1851 1072
rect -1783 1038 -1771 1072
rect -1863 1032 -1771 1038
rect -1705 1072 -1613 1078
rect -1705 1038 -1693 1072
rect -1625 1038 -1613 1072
rect -1705 1032 -1613 1038
rect -1547 1072 -1455 1078
rect -1547 1038 -1535 1072
rect -1467 1038 -1455 1072
rect -1547 1032 -1455 1038
rect -1389 1072 -1297 1078
rect -1389 1038 -1377 1072
rect -1309 1038 -1297 1072
rect -1389 1032 -1297 1038
rect -1231 1072 -1139 1078
rect -1231 1038 -1219 1072
rect -1151 1038 -1139 1072
rect -1231 1032 -1139 1038
rect -1073 1072 -981 1078
rect -1073 1038 -1061 1072
rect -993 1038 -981 1072
rect -1073 1032 -981 1038
rect -915 1072 -823 1078
rect -915 1038 -903 1072
rect -835 1038 -823 1072
rect -915 1032 -823 1038
rect -757 1072 -665 1078
rect -757 1038 -745 1072
rect -677 1038 -665 1072
rect -757 1032 -665 1038
rect -599 1072 -507 1078
rect -599 1038 -587 1072
rect -519 1038 -507 1072
rect -599 1032 -507 1038
rect -441 1072 -349 1078
rect -441 1038 -429 1072
rect -361 1038 -349 1072
rect -441 1032 -349 1038
rect -283 1072 -191 1078
rect -283 1038 -271 1072
rect -203 1038 -191 1072
rect -283 1032 -191 1038
rect -125 1072 -33 1078
rect -125 1038 -113 1072
rect -45 1038 -33 1072
rect -125 1032 -33 1038
rect 33 1072 125 1078
rect 33 1038 45 1072
rect 113 1038 125 1072
rect 33 1032 125 1038
rect 191 1072 283 1078
rect 191 1038 203 1072
rect 271 1038 283 1072
rect 191 1032 283 1038
rect 349 1072 441 1078
rect 349 1038 361 1072
rect 429 1038 441 1072
rect 349 1032 441 1038
rect 507 1072 599 1078
rect 507 1038 519 1072
rect 587 1038 599 1072
rect 507 1032 599 1038
rect 665 1072 757 1078
rect 665 1038 677 1072
rect 745 1038 757 1072
rect 665 1032 757 1038
rect 823 1072 915 1078
rect 823 1038 835 1072
rect 903 1038 915 1072
rect 823 1032 915 1038
rect 981 1072 1073 1078
rect 981 1038 993 1072
rect 1061 1038 1073 1072
rect 981 1032 1073 1038
rect 1139 1072 1231 1078
rect 1139 1038 1151 1072
rect 1219 1038 1231 1072
rect 1139 1032 1231 1038
rect 1297 1072 1389 1078
rect 1297 1038 1309 1072
rect 1377 1038 1389 1072
rect 1297 1032 1389 1038
rect 1455 1072 1547 1078
rect 1455 1038 1467 1072
rect 1535 1038 1547 1072
rect 1455 1032 1547 1038
rect 1613 1072 1705 1078
rect 1613 1038 1625 1072
rect 1693 1038 1705 1072
rect 1613 1032 1705 1038
rect 1771 1072 1863 1078
rect 1771 1038 1783 1072
rect 1851 1038 1863 1072
rect 1771 1032 1863 1038
rect 1929 1072 2021 1078
rect 1929 1038 1941 1072
rect 2009 1038 2021 1072
rect 1929 1032 2021 1038
rect 2087 1072 2179 1078
rect 2087 1038 2099 1072
rect 2167 1038 2179 1072
rect 2087 1032 2179 1038
rect 2245 1072 2337 1078
rect 2245 1038 2257 1072
rect 2325 1038 2337 1072
rect 2245 1032 2337 1038
rect -2235 971 -2189 983
rect -2235 181 -2229 971
rect -2195 181 -2189 971
rect -2235 169 -2189 181
rect -1919 971 -1873 983
rect -1919 181 -1913 971
rect -1879 181 -1873 971
rect -1919 169 -1873 181
rect -1603 971 -1557 983
rect -1603 181 -1597 971
rect -1563 181 -1557 971
rect -1603 169 -1557 181
rect -1287 971 -1241 983
rect -1287 181 -1281 971
rect -1247 181 -1241 971
rect -1287 169 -1241 181
rect -971 971 -925 983
rect -971 181 -965 971
rect -931 181 -925 971
rect -971 169 -925 181
rect -655 971 -609 983
rect -655 181 -649 971
rect -615 181 -609 971
rect -655 169 -609 181
rect -339 971 -293 983
rect -339 181 -333 971
rect -299 181 -293 971
rect -339 169 -293 181
rect -23 971 23 983
rect -23 181 -17 971
rect 17 181 23 971
rect -23 169 23 181
rect 293 971 339 983
rect 293 181 299 971
rect 333 181 339 971
rect 293 169 339 181
rect 609 971 655 983
rect 609 181 615 971
rect 649 181 655 971
rect 609 169 655 181
rect 925 971 971 983
rect 925 181 931 971
rect 965 181 971 971
rect 925 169 971 181
rect 1241 971 1287 983
rect 1241 181 1247 971
rect 1281 181 1287 971
rect 1241 169 1287 181
rect 1557 971 1603 983
rect 1557 181 1563 971
rect 1597 181 1603 971
rect 1557 169 1603 181
rect 1873 971 1919 983
rect 1873 181 1879 971
rect 1913 181 1919 971
rect 1873 169 1919 181
rect 2189 971 2235 983
rect 2189 181 2195 971
rect 2229 181 2235 971
rect 2189 169 2235 181
rect -2393 -181 -2347 -169
rect -2393 -971 -2387 -181
rect -2353 -971 -2347 -181
rect -2393 -983 -2347 -971
rect -2077 -181 -2031 -169
rect -2077 -971 -2071 -181
rect -2037 -971 -2031 -181
rect -2077 -983 -2031 -971
rect -1761 -181 -1715 -169
rect -1761 -971 -1755 -181
rect -1721 -971 -1715 -181
rect -1761 -983 -1715 -971
rect -1445 -181 -1399 -169
rect -1445 -971 -1439 -181
rect -1405 -971 -1399 -181
rect -1445 -983 -1399 -971
rect -1129 -181 -1083 -169
rect -1129 -971 -1123 -181
rect -1089 -971 -1083 -181
rect -1129 -983 -1083 -971
rect -813 -181 -767 -169
rect -813 -971 -807 -181
rect -773 -971 -767 -181
rect -813 -983 -767 -971
rect -497 -181 -451 -169
rect -497 -971 -491 -181
rect -457 -971 -451 -181
rect -497 -983 -451 -971
rect -181 -181 -135 -169
rect -181 -971 -175 -181
rect -141 -971 -135 -181
rect -181 -983 -135 -971
rect 135 -181 181 -169
rect 135 -971 141 -181
rect 175 -971 181 -181
rect 135 -983 181 -971
rect 451 -181 497 -169
rect 451 -971 457 -181
rect 491 -971 497 -181
rect 451 -983 497 -971
rect 767 -181 813 -169
rect 767 -971 773 -181
rect 807 -971 813 -181
rect 767 -983 813 -971
rect 1083 -181 1129 -169
rect 1083 -971 1089 -181
rect 1123 -971 1129 -181
rect 1083 -983 1129 -971
rect 1399 -181 1445 -169
rect 1399 -971 1405 -181
rect 1439 -971 1445 -181
rect 1399 -983 1445 -971
rect 1715 -181 1761 -169
rect 1715 -971 1721 -181
rect 1755 -971 1761 -181
rect 1715 -983 1761 -971
rect 2031 -181 2077 -169
rect 2031 -971 2037 -181
rect 2071 -971 2077 -181
rect 2031 -983 2077 -971
rect 2347 -181 2393 -169
rect 2347 -971 2353 -181
rect 2387 -971 2393 -181
rect 2347 -983 2393 -971
rect -2337 -1038 -2245 -1032
rect -2337 -1072 -2325 -1038
rect -2257 -1072 -2245 -1038
rect -2337 -1078 -2245 -1072
rect -2179 -1038 -2087 -1032
rect -2179 -1072 -2167 -1038
rect -2099 -1072 -2087 -1038
rect -2179 -1078 -2087 -1072
rect -2021 -1038 -1929 -1032
rect -2021 -1072 -2009 -1038
rect -1941 -1072 -1929 -1038
rect -2021 -1078 -1929 -1072
rect -1863 -1038 -1771 -1032
rect -1863 -1072 -1851 -1038
rect -1783 -1072 -1771 -1038
rect -1863 -1078 -1771 -1072
rect -1705 -1038 -1613 -1032
rect -1705 -1072 -1693 -1038
rect -1625 -1072 -1613 -1038
rect -1705 -1078 -1613 -1072
rect -1547 -1038 -1455 -1032
rect -1547 -1072 -1535 -1038
rect -1467 -1072 -1455 -1038
rect -1547 -1078 -1455 -1072
rect -1389 -1038 -1297 -1032
rect -1389 -1072 -1377 -1038
rect -1309 -1072 -1297 -1038
rect -1389 -1078 -1297 -1072
rect -1231 -1038 -1139 -1032
rect -1231 -1072 -1219 -1038
rect -1151 -1072 -1139 -1038
rect -1231 -1078 -1139 -1072
rect -1073 -1038 -981 -1032
rect -1073 -1072 -1061 -1038
rect -993 -1072 -981 -1038
rect -1073 -1078 -981 -1072
rect -915 -1038 -823 -1032
rect -915 -1072 -903 -1038
rect -835 -1072 -823 -1038
rect -915 -1078 -823 -1072
rect -757 -1038 -665 -1032
rect -757 -1072 -745 -1038
rect -677 -1072 -665 -1038
rect -757 -1078 -665 -1072
rect -599 -1038 -507 -1032
rect -599 -1072 -587 -1038
rect -519 -1072 -507 -1038
rect -599 -1078 -507 -1072
rect -441 -1038 -349 -1032
rect -441 -1072 -429 -1038
rect -361 -1072 -349 -1038
rect -441 -1078 -349 -1072
rect -283 -1038 -191 -1032
rect -283 -1072 -271 -1038
rect -203 -1072 -191 -1038
rect -283 -1078 -191 -1072
rect -125 -1038 -33 -1032
rect -125 -1072 -113 -1038
rect -45 -1072 -33 -1038
rect -125 -1078 -33 -1072
rect 33 -1038 125 -1032
rect 33 -1072 45 -1038
rect 113 -1072 125 -1038
rect 33 -1078 125 -1072
rect 191 -1038 283 -1032
rect 191 -1072 203 -1038
rect 271 -1072 283 -1038
rect 191 -1078 283 -1072
rect 349 -1038 441 -1032
rect 349 -1072 361 -1038
rect 429 -1072 441 -1038
rect 349 -1078 441 -1072
rect 507 -1038 599 -1032
rect 507 -1072 519 -1038
rect 587 -1072 599 -1038
rect 507 -1078 599 -1072
rect 665 -1038 757 -1032
rect 665 -1072 677 -1038
rect 745 -1072 757 -1038
rect 665 -1078 757 -1072
rect 823 -1038 915 -1032
rect 823 -1072 835 -1038
rect 903 -1072 915 -1038
rect 823 -1078 915 -1072
rect 981 -1038 1073 -1032
rect 981 -1072 993 -1038
rect 1061 -1072 1073 -1038
rect 981 -1078 1073 -1072
rect 1139 -1038 1231 -1032
rect 1139 -1072 1151 -1038
rect 1219 -1072 1231 -1038
rect 1139 -1078 1231 -1072
rect 1297 -1038 1389 -1032
rect 1297 -1072 1309 -1038
rect 1377 -1072 1389 -1038
rect 1297 -1078 1389 -1072
rect 1455 -1038 1547 -1032
rect 1455 -1072 1467 -1038
rect 1535 -1072 1547 -1038
rect 1455 -1078 1547 -1072
rect 1613 -1038 1705 -1032
rect 1613 -1072 1625 -1038
rect 1693 -1072 1705 -1038
rect 1613 -1078 1705 -1072
rect 1771 -1038 1863 -1032
rect 1771 -1072 1783 -1038
rect 1851 -1072 1863 -1038
rect 1771 -1078 1863 -1072
rect 1929 -1038 2021 -1032
rect 1929 -1072 1941 -1038
rect 2009 -1072 2021 -1038
rect 1929 -1078 2021 -1072
rect 2087 -1038 2179 -1032
rect 2087 -1072 2099 -1038
rect 2167 -1072 2179 -1038
rect 2087 -1078 2179 -1072
rect 2245 -1038 2337 -1032
rect 2245 -1072 2257 -1038
rect 2325 -1072 2337 -1038
rect 2245 -1078 2337 -1072
rect -136 -1176 136 -1170
rect -136 -1210 -124 -1176
rect 124 -1210 136 -1176
rect -136 -1216 136 -1210
<< properties >>
string FIXED_BBOX -2504 -1193 2504 1193
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 10.0 l 0.5 m 1 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 5 viagr 0 viagl 0 viagt 0
<< end >>
